#Version=1.16
#Author= Hans Eriksson, E-mail: hans.ericson@bredband.net
reversed = (omv�nd f�rg)
A00.7=Anderssens �ppning
A00.8=Hemsk krypande (Basmans) �ppning 
A00.6=Wares (h�-�ngs) �ppning
A00.11=Durkins attack
A00.18=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning
A00.19=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...Nf6
A00.20=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...Nf6 2.Nf3
A00.21=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: T�bingen gambit
A00.22=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...e5
A00.23=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...e5 2.Nf3
A00.24=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: Sicilianska varianten
A00.25=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: Sicilianska varianten, 2.Nf3
A00.26=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: Sicilianska varianten, 2.Nf3 Nc6
A00.27=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5
A00.28=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5 2.Nf3
A00.29=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5 2.Nf3 Nf6
A00.30=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5 2.e4
A00.31=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5 2.e4 d4
A00.32=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: 1...d5 2.e4 dxe4
A00.33=Dunsts (Sleipner-Heinrichsen-Van Geet) �ppning: Hectors gambit
A00.46=Polsk (Sokolsky-Orangutang) �ppning
A00.47=Polsk (Sokolsky-Orangutang) �ppning: Birminghams gambit
A00.48=Polsk (Sokolsky-Orangutang) �ppning: 1...Nf6
A00.49=Polsk (Sokolsky-Orangutang) �ppning: 1...Nf6 2.Bb2
A00.50=Polsk (Sokolsky-Orangutang) �ppning: Gligoric-Smyslovvarianten, 1...Nf6 2.Bb2 e6
A00.51=Polsk (Sokolsky-Orangutang) �ppning: Utflankeringsvarianten, 1...c6
A00.52=Polsk (Sokolsky-Orangutang) �ppning: Sch�hlers gambit
A00.53=Polsk (Sokolsky-Orangutang) �ppning: 1...d5
A00.54=Polsk (Sokolsky-Orangutang) �ppning: 1...d5 2.Bb2
A00.55=Polsk (Sokolsky-Orangutang) �ppning: 1...d5 2.Bb2 Bf5
A00.56=Polsk (Sokolsky-Orangutang) �ppning: Golombeksvarianten
A00.57=Polsk (Sokolsky-Orangutang) �ppning: Golombeksvarianten, 1...d5 2.Bb2 Nf6 3.e3
A00.58=Polsk (Sokolsky-Orangutang) �ppning: 1...e5
A00.59=Polsk (Sokolsky-Orangutang) �ppning: Bugayevattacken
A00.60=Polsk (Sokolsky-Orangutang) �ppning: 1...e5 2.Bb2
A00.61=Polsk (Sokolsky-Orangutang) �ppning: Wolfertz gambit
A00.64=Polsk (Sokolsky-Orangutang) �ppning: Taimanovarianten, 1...e5 2.Bb2 d6
A00.62=Polsk (Sokolsky-Orangutang) �ppning: 1...e5 2.Bb2 f6
A00.63=Polsk (Sokolsky-Orangutang) �ppning: Schiffler-Tartakower gambit
A00.65=Polsk (Sokolsky-Orangutang) �ppning: Avbytesvarianten, 2...Bxb4
A00.66=Polsk (Sokolsky-Orangutang) �ppning: Avbytesvarianten, 2...Bxb4 3.Bxe5
A00.67=Polsk (Sokolsky-Orangutang) �ppning: Avbytesvarianten, 2...Bxb4 3.Bxe5 Nf6
A00.68=Polsk (Sokolsky-Orangutang) �ppning: Avbytesvarianten, 2...Bxb4 3.Bxe5 Nf6 4.c4
A00.69=Polsk (Sokolsky-Orangutang) �ppning: Avbytesvarianten, 2...Bxb4 3.Bxe5 Nf6 4.Nf3
A00.12=Saragossas �ppning
A00.13=Mieses �ppning
A00.15=Mieses �ppning: 1...d5
A00.14=Mieses �ppning: 1...e5
A00.16=Avb�jd tagg�ppning
A00.17=Van Kruijs �ppning
A00.2=Barnes (T�lamods) �ppning
A00.3=Hammerschlags (Stekt r�v-fl�skkotlett) �ppning
A00.9=Amars (Paris) �ppning
A00.10=Amars (Paris) �ppning: Paris gambit
A00.70=Benkos �ppning
A00.74=Benkos �ppning: 1...d5
A00.75=Benkos �ppning: 1.g3 d5 2.Bg2
A00.76=Benkos �ppning: 1.g3 d5 2.Bg2 c6
A00.77=Benkos �ppning: 1.g3 d5 2.Bg2 e5
A00.78=Benkos �ppning: 1.g3 d5 2.Bg2 Nf6
A00.73=Benkos �ppning: Reti-Antagen Kungsindisk-Engelsk transposition, 1...e5
A00.72=Benkos �ppning: Symmetrisk
A00.71=Benkos �ppning: 1...Nf6
A00.34=Grobs (Fric-Kilibr) �ppning
A00.35=Grobs (Fric-Kilibr) �ppning: Alessis gambit
A00.36=Grobs (Fric-Kilibr) �ppning: Dubbel Grob
A00.37=Grobs (Fric-Kilibr) �ppning: 1...e5
A00.38=Grobs (Fric-Kilibr) �ppning: 1...d5
A00.39=Grobs gambit
A00.40=Grobs gambit: 2...e5
A00.41=Grobs gambit: Hurstattacken
A00.42=Grobs gambit: 2...c6
A00.43=Grobs gambit: Taggattacken
A00.44=Antagen Grobs gambit
A00.45=Antagen Grobs gambit: Fritz gambit
A00.5=Clemenz (Mead-Basman-de Klerk-Welling) �ppning
A00.4=Kadas (Desprez) �ppning
A01.1=Nimzowitsch-Larsen attack
A01.2=Nimzowitsch-Larsen attack: Polsk variant
A01.3=Nimzowitsch-Larsen attack: Symmetrisk variant
A01.4=Nimzowitsch-Larsen attack: Holl�ndsk variant
A01.5=Nimzowitsch-Larsen attack: Ringelbachs gambit
A01.6=Nimzowitsch-Larsen attack: Engelska varianten
A01.7=Nimzowitsch-Larsen attack: Indiska varianten
A01.8=Nimzowitsch-Larsen attack: Indiska varianten, 1.b3 Nf6 2.Bb2 g6
A01.9=Nimzowitsch-Larsen attack: Taggvarianten
A01.10=Nimzowitsch-Larsen attack: Klassiska varianten, 1...d5
A01.11=Nimzowitsch-Larsen attack: Klassiska varianten, 1...d5 2.Bb2
A01.12=Nimzowitsch-Larsen attack: Moderna varianten, 1...e5
A01.13=Nimzowitsch-Larsen attack: Moderna varianten, 1...e5 2.Bb2
A01.14=Nimzowitsch-Larsen attack: Moderna varianten, 1...e5 2.Bb2 d6
A01.15=Nimzowitsch-Larsen attack: Moderna varianten, 1...e5 2.Bb2 Nc6
A01.16=Nimzowitsch-Larsen attack: Moderna varianten, Paschmanns gambit
A01.17=Nimzowitsch-Larsen attack: Moderna varianten, 1...e5 2.Bb2 Nc6 3.e3
A02.1=Birds �ppning
A02.2=Birds �ppning: Hobbs gambit
A02.3=Birds �ppning: Symmetriska varianten
A02.4=Birds �ppning: Schweizisk gambit
A02.5=Birds �ppning: Antagen Schweizisk gambit
A02.6=Birds �ppning: 1..d6
A02.7=Birds �ppning: 1..g6
A02.8=Birds �ppning: 1.f4 g6 2.Nf3 Bg7 3.e3
A02.9=Birds �ppning: 1.f4 g6 2.Nf3 Bg7 3.g3
A02.10=Birds �ppning: 1..c5
A02.11=Birds �ppning: 1..c5 2.Nf3 Nc6
A02.12=Birds �ppning: Froms gambit
A02.13=Birds �ppning: Froms gambit Antagen
A02.14=Birds �ppning: Froms gambit, Schlecter
A02.15=Birds �ppning: Froms gambit, 2...d6
A02.16=Birds �ppning: Froms gambit, 3.exd6
A02.17=Birds �ppning: Froms gambit, Langheld gambit
A02.18=Birds �ppning: Froms gambit, 3...Bxd6
A02.19=Birds �ppning: Froms gambit, Lipke
A02.20=Birds �ppning: Froms gambit, Laskervarianten
A02.21=Birds �ppning: Froms gambit, Lasker, 5.d4
A02.22=Birds �ppning: Froms gambit, Lasker, Dambytevarianten
A02.23=Birds �ppning: Froms gambit, Lasker, 5.g3
A02.24=Birds �ppning: 1..Nf6
A02.25=Birds �ppning: 1..Nf6 2.g3
A02.26=Birds �ppning: 1..Nf6 2.e3
A02.27=Birds �ppning: 1..Nf6 2.b3
A02.28=Birds �ppning: 1..Nf6 2.Nf3
A02.29=Birds �ppning: 1..Nf6 2.Nf3 d6
A02.30=Birds �ppning: 1..Nf6 2.Nf3 c5
A02.31=Birds �ppning: 1..Nf6 2.Nf3 g6
A02.32=Birds �ppning: Batavo Polsk attack
A02.33=Birds �ppning: 1..Nf6 2.Nf3 g6 3.g3
A02.34=Birds �ppning: Mortars attack 1.. Nf6 2.Nf3 g6 3.g3 Bg7 4.Bg2
A02.35=Birds �ppning: Mortars attack, 4.Bg2 d6
A03.1=Birds �ppning: 1...d5
A03.2=Birds �ppning: Dudweilers gambit
A03.3=Birds �ppning: Mujannah-Sturms gambit
A03.4=Birds �ppning: Williams gambit
A03.5=Birds �ppning: 1.f4 d5 2.b3
A03.6=Birds �ppning: 1.f4 d5 2.b3 Nf6
A03.7=Birds �ppning: 1.f4 d5 2.b3 Nf6 3.Bb2
A03.8=Birds �ppning: 1.f4 d5 2.g3
A03.9=Birds �ppning: 1.f4 d5 2.g3 Nf6
A03.10=Birds �ppning: 1.f4 d5 2.g3 Nf6 3.Bg2
A03.11=Birds �ppning: Laskervarianten
A03.12=Birds �ppning: Laskervarianten
A03.13=Birds �ppning: 1...d5 2.Nf3
A03.14=Birds �ppning: 1...d5 2.Nf3 c5
A03.15=Birds �ppning: Batavos gambit
A03.16=Birds �ppning: 1...d5 2.Nf3 c5 3.e3
A03.17=Birds �ppning: 1...d5 2.Nf3 g6
A03.18=Birds �ppning: 1...d5 2.Nf3 g6 3.e3
A03.19=Birds �ppning: 1...d5 2.Nf3 g6 3.g3
A03.20=Birds �ppning: 1...d5 2.Nf3 g6 3.g3 Bg7 4.Bg2
A03.21=Birds �ppning: 1...d5 2.Nf3 Nf6
A03.22=Birds �ppning: 1...d5 2.Nf3 Nf6 3.b3
A03.23=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3
A03.24=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6
A03.25=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6 4.Bg2 Bg7
A03.26=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6 4.Bg2 Bg7 5.d3
A03.27=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6: 5.O-O
A03.28=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6: 5.O-O O-O
A03.29=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6: 5.O-O O-O 6.d3
A03.30=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6: 6.d3 c6
A03.31=Birds �ppning: 1...d5 2.Nf3 Nf6 3.g3 g6: 6.d3 c5
A03.32=Birds �ppning: Laskervarianten
A03.33=Birds �ppning: Laskervarianten, 3...Bg4
A03.34=Birds �ppning: Laskervarianten, 3...e6
A03.35=Birds �ppning: Laskervarianten, 3...c5
A03.36=Birds �ppning: Laskervarianten, 3...c5 4.b3
A03.37=Birds �ppning: Laskervarianten, 3...g6
A04.1=Retis �ppning
A04.2=Retis �ppning: Herrstr�ms gambit
A04.3=Retis �ppning: 1...b6
A04.4=Retis �ppning: 1...b5
A04.5=Retis �ppning: 1...Nc6
A04.6=Retis �ppning: 1...e6
A04.7=Retis �ppning: 1...e6 2.g3
A04.8=Retis �ppning: 1...g6
A04.9=Retis �ppning: 1...g6 2.g3
A04.10=Retis �ppning: 1...g6 2.g3 Bg7
A04.11=Retis �ppning: 1...g6 2.g3 Bg7 3.Bg2
A04.12=Retis �ppning: 1...f5
A04.13=Retis �ppning: 1...f5 2.d3
A04.14=Retis �ppning: 1...f5 2.d3 Nf6
A04.15=Retis �ppning: Avb�jd Lisitsins gambit
A04.16=Retis �ppning: 1...f5 2.g3
A04.17=Retis �ppning: Lisitsins gambit
A04.18=Retis �ppning: Lisitsins gambit: 3.Ng5 Nf6
A04.19=Retis �ppning: Lisitsins gambit: 3.Ng5 Nf6 4.d3 e5
A04.20=Retis �ppning: Lisitsins gambit: 3.Ng5 Nf6 4.d3 e3
A04.21=Retis �ppning: Lisitsins gambit: 3.Ng5 e5
A04.22=Retis �ppning: Lisitsins gambit: 3.Ng5 d5
A04.23=Retis �ppning: 1...d6
A04.24=Retis �ppning: 1...c5
A04.25=Retis �ppning: 1...c5, Nimzowitsch-Larsen
A04.26=Retis �ppning: 1...c5 2.g3
A04.27=Retis �ppning: 1...c5 2.g3 b6
A04.28=Retis �ppning: 1...c5 2.g3 b6 3.Bg2 Bb7
A04.29=Retis �ppning: 1...c5 2.g3 g6
A04.30=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7
A04.31=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6
A04.32=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6 5.d3
A04.33=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6 5.d3 Nf6 6.e4
A04.34=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6 5.d3 Nf6
A04.35=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6 5.d3 d6 6.e4
A04.36=Retis �ppning: 1...c5 2.g3 g6 3.Bg2 Bg7 4.O-O Nc6 5.d3 e6 6.e4
A04.37=Retis �ppning: 1...c5 2.g3 Nc6
A04.38=Retis �ppning: 1...c5 2.g3 Nc6 3.Bg2
A05.1=Retis �ppning: 1...Nf6
A05.2=Retis �ppning: 1...Nf6 2.b3
A05.3=Retis �ppning: Santasieres Folly
A05.4=Retis �ppning: 1...Nf6 2.e3
A05.5=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3
A05.6=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 c5
A05.7=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 c5 3.Bg2
A05.8=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 c5 3.Bg2 Nc6
A05.9=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 b6
A05.10=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 b6 3.Bg2
A05.11=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 b6 3.Bg2 Bb7
A05.12=Retis �ppning: Antagen Kungsindisk, Spasskyvarianten 1.Nf3 Nf6 2.g3 b5
A05.13=Retis �ppning: Antagen Kungsindisk, Spasskyvarianten 1.Nf3 Nf6 2.g3 b5 3.Bg2
A05.14=Retis �ppning: Antagen Kungsindisk, 1.Nf3 Nf6 2.g3 g6
A05.15=Retis �ppning: Antagen Kungsindisk, Reti-Smyslovvarianten 3.b4
A05.16=Retis �ppning: Antagen Kungsindisk, Reti-Smyslovvarianten 3.b4 Bg7 5.Bb2
A05.17=Retis �ppning: Antagen Kungsindisk, 3.Bg2
A05.18=Retis �ppning: Antagen Kungsindisk, 3.Bg2 Bg7
A05.19=Retis �ppning: Antagen Kungsindisk, 3.Bg2 Bg7 4.O-O
A05.20=Retis �ppning: Antagen Kungsindisk, 3.Bg2 Bg7 4.O-O O-O
A05.21=Retis �ppning: Antagen Kungsindisk, 3.Bg2 Bg7 4.O-O O-O 5.d3
A05.23=Retis �ppning: Antagen Kungsindisk, 3.Bg2 Bg7 4.O-O O-O 5.d3 d6
A06.1=Retis �ppning: 1...d5
A06.2=Retis �ppning: Gammaindisk attack
A06.3=Retis �ppning: Gammalindisk attack, 1.Nf3 d5 2.d3 Nf6
A06.4=Retis �ppning: 1...d5 2.e3
A06.5=Retis �ppning: Santasieres Folly, 1.Nf3 d5 2.b4
A06.6=Retis �ppning: Santasieres Folly, 1.Nf3 d5 2.b4 Nf6
A06.7=Retis �ppning: Tennisons (Zukertort-Lemberg) gambit
A06.8=Retis �ppning: Antagen Tennisons (Zukertort-Lemberg) gambit
A06.9=Retis �ppning: Nimzowitsch-Larsen
A06.10=Retis �ppning: Nimzowitsch-Larsen, 2...c5
A06.11=Retis �ppning: Nimzowitsch-Larsen, 2...Bg4
A06.12=Retis �ppning: Nimzowitsch-Larsen, 2...Bg4 3.Bb2
A06.13=Retis �ppning: Nimzowitsch-Larsen, 2...Bg43.Bb2 Nd7 4.e3
A06.14=Retis �ppning: Nimzowitsch-Larsen, 2...Nf6
A06.15=Retis �ppning: Nimzowitsch-Larsen, 2...Nf6 3.Bb2
A06.16=Retis �ppning: Nimzowitsch-Larsen, 2...Nf6 Nf6 3.Bb2 e6
A06.17=Retis �ppning: Nimzowitsch-Larsen, 2...Nf6 Nf6 3.Bb2 e6 4.e3
A07.1=Retis �ppning: Antagen Kungsindisk, 2.g3
A07.2=Retis �ppning: Antagen Kungsindisk, 2.g3 Nc6
A07.3=Retis �ppning: Antagen Kungsindisk, 2.g3 Nc6 3.Bg2 e5
A07.4=Retis �ppning: Antagen Kungsindisk, 2.g3 Nc6 3.Bg2 e5 4.d3 Nf6
A07.5=Retis �ppning: Antagen Kungsindisk, 2.g3 Nc6 3.Bg2 e5 4.d3 Nf6 5.O-O
A07.6=Retis �ppning: Antagen Kungsindisk, 2.g3 Nc6 3.Bg2 e5 4.d3 Nf6 5.O-O Be7
A07.7=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten
A07.8=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 Bg4
A07.9=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 Bg4 4.O-O
A07.10=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 Bg4 4.O-O Nd7
A07.11=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 Bg4 4.O-O Nd7 5.d3
A07.12=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 c6 4.O-O Bg4
A07.13=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, 3.Bg2 c6 4.O-O Bg4 5.d3
A07.14=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, Huvudvarianten
A07.15=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, Huvudvarianten, 6.Nbd2
A07.16=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, Huvudvarianten, 6.Nbd2 e6
A07.17=Retis �ppning: Antagen Kungsindisk, Jugoslaviska varianten, Huvudvarianten, 6.Nbd2 e5
A07.18=Retis �ppning: Antagen Kungsindisk, Keresvarianten
A07.19=Retis �ppning: Antagen Kungsindisk, Keresvarianten, 3.Bg2 Nd7
A07.20=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 Nf6
A07.21=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 Nf6 3.Bg2
A07.22=Retis �ppning: Antagen Kungsindisk, Neo-Gr�nfeldvarianten
A07.23=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 Nf6 3.Bg2 Bf5
A07.24=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 Nf6 3.Bg2 e6
A07.25=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 Nf6 3.Bg2 c6
A07.26=Retis �ppning: Antagen Kungsindisk, Petrosianvarianten
A07.27=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 g6
A07.28=Retis �ppning: Antagen Kungsindisk, 1.Nf3 d5 2.g3 g6 3.Bg2
A07.29=Retis �ppning: Antagen Kungsindisk, Pachmanssystemet, 3...Bg7 4.O-O e5 5.d3 Ne7
A08.1=Retis �ppning: Antagen Kungsindisk, 2...c5
A08.2=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2
A08.3=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 g6 4.O-O Bg7
A08.4=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 g6 4.O-O Bg7 5.d3
A08.5=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 g6 4.O-O Bg7 5.d3 Nf6
A08.6=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 g6 4.O-O Bg7 5.d3 Nf6 6.Nbd2 O-O
A08.7=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 g6 4.O-O Nc6 5.d3 Nf6
A08.8=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 Nc6
A08.9=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 Nc6 4.O-O
A08.11=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 Nf6
A08.12=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 Nf6 4.O-O
A08.13=Retis �ppning: Antagen Kungsindisk, 2...c5 3.Bg2 Nf6 4.O-O Nc6
A08.14=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nge7 6.Nbd2 b6 7.e4
A08.15=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nf6 6.Nbd2 b6 7.e4
A08.16=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nge7 6.Nbd2 g6 7.e4 Bg7
A08.17=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nf6 6.Nbd2 g6 7.e4 Bg7
A08.18=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nf6 6.Nbd2 Be7 7.e4
A08.19=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Nf6 6.Nbd2 Be7 7.e4 O-O 8.Re1
A08.20=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Bd6 6.Nbd2 Nge7 7.e4
A08.21=Retis �ppning: Antagen Kungsindisk, Fransk, 3...Nc6 4.O-O e6 5.d3 Bd6 6.Nbd2 Nge7 7.e4 O-O 8.Re1
A09.1=Retis �ppning: 2.c4
A09.2=Retis �ppning: Avanceravarianten
A09.3=Retis �ppning: Avanceravarianten, Engelsk-Polsk attack
A09.4=Retis �ppning: Avanceravarianten, Engelsk-Polsk attack, 3...g6
A09.5=Retis �ppning: Avanceravarianten, 3.e3
A09.6=Retis �ppning: Avanceravarianten, 3.e3 c5
A09.7=Retis �ppning: Avanceravarianten, 3.e3 Nc6
A09.8=Retis �ppning: Avanceravarianten, 3.e3 Nc6 4.exd4 Nxd4
A09.9=Retis �ppning: Avanceravarianten, 3.g3
A09.10=Retis �ppning: Avanceravarianten, 3.g3 Nc6
A09.11=Retis �ppning: Avanceravarianten, 3.g3 Nc6 4.Bg2 e5
A09.12=Retis �ppning: Avanceravarianten, 3.g3 g6
A09.13=Retis �ppning: Avanceravarianten, 3.g3 g6 4.Bg2 Bg7
A09.14=Retis �ppning: Avanceravarianten, 3.g3 c5
A09.15=Retis �ppning: Avanceravarianten, 3.g3 c5 4.Bg2 Nc6
A09.16=Retis �ppning: Avanceravarianten, 3.g3 c5 4.Bg2 Nc6 5.d3 e5
A09.17=Retis �ppning: Antagen
A09.18=Retis �ppning: Antagen, 3.g3
A09.19=Retis �ppning: Antagen, 3.g3 e6
A09.20=Retis �ppning: Antagen, 3.Qa4+
A09.21=Retis �ppning: Antagen, 3.Na3
A09.22=Retis �ppning: Antagen, 3.Na3 a6
A09.23=Retis �ppning: Antagen, 3.Na3 c5
A09.24=Retis �ppning: Antagen, 3.e3
A09.25=Retis �ppning: Antagen, Keresvarianten
A09.26=Retis �ppning: Antagen, 3.e3 Nf6
A09.27=Retis �ppning: Antagen, 3.e3 Nf6 4.Bxc4 e6
A10.1=Engelskt
A10.2=Engelskt: 1...g5
A10.3=Engelskt: 1...g5 2.d4
A10.4=Engelskt: Myers gambit
A10.5=Engelskt: 1...Nc6
A10.6=Engelskt: 1...Nc6 2.Nc3
A10.7=Engelskt: J�nisch gambit
A10.8=Engelskt: Vector
A10.9=Engelskt: 1...b6
A10.10=Engelskt: 1...b6 2.Nf3
A10.11=Engelskt: 1...b6 2.Nf3 Bb7
A10.12=Engelskt: 1...b6 2.Nc3
A10.13=Engelskt: 1...b6 2.Nc3 e6
A10.14=Engelskt: 1...b6 2.Nc3 e6 3.e4
A10.15=Engelskt: 1...b6 2.Nc3 Bb7
A10.16=Engelskt: 1...b6 2.Nc3 Bb7 3.e4
A10.17=Engelskt: 1...b6 2.Nc3 Bb7 3.e4 e6
A10.18=Engelskt: 1...d6
A10.19=Engelskt: 1...d6 2.Nc3
A10.20=Engelskt: 1...d6 2.Nf3
A10.21=Engelskt: 1...g6
A10.22=Engelskt: 1...g6 2.g3
A10.23=Engelskt: 1...g6 2.Nc3
A10.24=Engelskt: 1...g6 2.Nc3 Bg7
A10.25=Engelskt: 1...g6 2.Nc3 Bg7 3.g3
A10.26=Engelskt: 1...g6 2.Nf3
A10.27=Engelskt: 1...g6 2.Nf3 Bg7
A10.28=Engelskt: 1...g6 2.e4
A10.29=Engelskt: Adorjan f�rsvar
A10.30=Engelskt: Engelsk-Holl�ndsk
A10.31=Engelskt: Wades gambit
A10.32=Engelskt: Engelsk-Holl�ndsk, 2.g3
A10.33=Engelskt: Engelsk-Holl�ndsk, 2.g3 Nf6
A10.34=Engelskt: Engelsk-Holl�ndsk, 2.g3 Nf6 3.Bg2
A10.35=Engelskt: Engelsk-Holl�ndsk, 2.Nc3
A10.36=Engelskt: Engelsk-Holl�ndsk, 2.Nc3 Nf6
A10.37=Engelskt: Engelsk-Holl�ndsk, 2.Nc3 Nf6 3.g3
A10.38=Engelskt: Engelsk-Holl�ndsk, 2.Nc3 Nf6 3.g3 g6
A10.39=Engelskt: Engelsk-Holl�ndsk, 2.Nf3
A10.40=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 e6
A10.41=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6
A10.42=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.Nc3
A10.43=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3
A10.44=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6
A10.45=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2
A10.46=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2 c6 5.O-O d5
A10.47=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2 Be7
A10.48=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2 Be7 5.O-O
A10.49=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2 Be7 5.O-O O-O
A10.50=Engelskt: Engelsk-Holl�ndsk, 2.Nf3 Nf6 3.g3 e6 4.Bg2 Be7 5.O-O O-O 6.Nc3
A11.1=Engelskt: Caro-Kann f�rsvar
A11.2=Engelskt: Caro-Kann f�rsvar, 2.g3
A11.3=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6
A11.4=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5
A11.5=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3
A11.6=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3 Bf5
A11.7=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3 Bf5 5.O-O
A11.8=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3 Bf5 5.O-O e6 6.d3
A11.9=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3 Bg4
A11.10=Engelskt: Caro-Kann f�rsvar, 2.g3 Nf6 3.Bg2 d5 4.Nf3 Bg4 5.O-O
A11.11=Engelskt: Caro-Kann f�rsvar, 2.Nc3
A11.12=Engelskt: Caro-Kann f�rsvar, 2.Nc3 d5
A11.13=Engelskt: Caro-Kann f�rsvar, 2.Nf3
A11.14=Engelskt: Caro-Kann f�rsvar, 2.Nf3 Nf6
A11.15=Engelskt: Caro-Kann f�rsvar, 2.Nf3 d5
A11.16=Engelskt: Caro-Kann f�rsvar, 3.g3
A11.17=Engelskt: Caro-Kann f�rsvar, 3.g3 Bg4
A11.18=Engelskt: Caro-Kann f�rsvar, 3.g3 Bg4 4.Bg2
A11.19=Engelskt: Caro-Kann f�rsvar, 3.e3
A11.20=Engelskt: Caro-Kann f�rsvar, 3.e3 Nf6
A11.21=Engelskt: Caro-Kann f�rsvar, 3.e3 Nf6 4.Nc3
A12.1=Engelskt: Caro-Kann f�rsvar, 3.b3
A12.2=Engelskt: Torref�rsvar, 3.b3 Nf6 4.g3 Bg4
A12.3=Engelskt: Torref�rsvar, 3.b3 Nf6 4.g3 Bg4 5.Bg2
A12.4=Engelskt: Torref�rsvar, 3.b3 Nf6 4.g3 Bg4 5.Bg2 e6
A12.5=Engelskt: Torref�rsvar, 3.b3 Nf6 4.g3 Bg4 5.Bg2 e6 6.Bb2
A12.6=Engelskt: Londonf�rsvar, 4...Bf5
A12.7=Engelskt: Londonf�rsvar, 4...Bf5 5.Bg2
A12.8=Engelskt: Londonf�rsvar, 4...Bf5 5.Bg2 e6
A12.9=Engelskt: Londonf�rsvar, 4...Bf5 5.Bg2 e6 6.Bb2
A12.10=Engelskt: Caro-Kannf�rsvar, 3.b3 Nf6 4.Bb2
A12.11=Engelskt: Bledvarianten, 4...g6
A12.12=Engelskt: Bledvarianten, 4...g6 5.e3 Bg7
A12.13=Engelskt: New York-London f�rsvaret
A12.14=Engelskt: Capablancavarianten
A12.15=Engelskt: Bogoljubowvarianten
A13.1=Engelskt: 1...e6
A13.2=Engelskt: 1...e6 2.g3
A13.3=Engelskt: 1...e6 2.g3 d5
A13.4=Engelskt: 1...e6 2.g3 d5
A13.5=Engelskt: 1...e6 2.Nc3
A13.6=Engelskt: 1...e6 2.Nc3 Bb4
A13.7=Engelskt: 1...e6 2.Nc3 d5
A13.8=Engelskt: 1...e6 2.Nf3
A13.9=Engelskt: 1...e6 2.Nf3 Nf6
A13.10=Engelskt: 1...e6 2.Nf3 Nf6 3.g3
A13.11=Engelskt: Romanishins gambit
A13.12=Engelskt: 1...e6 2.Nf3 d5
A13.13=Engelskt: Agincourtvarianten,  3.b3
A13.14=Engelskt: Wimpeysystemet, 3.b3 Nf6 4.Bb2 c5 5.e3
A13.15=Engelskt: Wimpeysystemet, 3.b3 Nf6 4.Bb2 c5 5.e3 Nc6
A13.16=Engelskt: Agincourtvarianten, 3.g3
A13.17=Engelskt: Kurajicas f�rsvar
A13.18=Engelskt: Kurajicas f�rsvar,  4.Qc2
A13.19=Engelskt: Neo-Katalansk
A13.20=Engelskt: Neo-Katalansk, 4.Bg2
A13.21=Engelskt: Neo-Katalansk, 4...c6
A13.22=Engelskt: Neo-Katalansk, 4...c6 5.b3
A13.23=Engelskt: Neo-Katalansk, 4...c5
A13.24=Engelskt: Neo-Katalansk, 4...c5 5.O-O
A13.25=Engelskt: Antagen Neo-Katalansk
A13.26=Engelskt: Antagen Neo-Katalansk, 5.Qa4+
A13.27=Engelskt: Antagen Neo-Katalansk, 5.Qa4+ Nbd7
A13.28=Engelskt: Antagen Neo-Katalansk, 5.Qa4+ Nbd7 6.O-O
A13.29=Engelskt: Antagen Neo-Katalansk, 5.Qa4+ Nbd7 6.Qxc4
A13.30=Engelskt: Antagen Neo-Katalansk, 5.Qa4+ Nbd7 6.Qxc4 a6
A13.31=Engelskt: Antagen Neo-Katalansk, 5.Qa4+ Nbd7 6.Qxc4 c5
A14.1=Engelskt: Avb�jd Neo-Katalansk
A14.2=Engelskt: Avb�jd Neo-Katalansk
A14.3=Engelskt: Avb�jd Neo-Katalansk, 5...c6
A14.4=Engelskt: Avb�jd Neo-Katalansk, 5...c5
A14.5=Engelskt: Avb�jd Neo-Katalansk, 5...O-O
A14.6=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3
A14.7=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 b6
A14.8=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 b6 7.Bb2 Bb7
A14.9=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 b6 7.Bb2 Bb7 8.e3
A14.10=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 c5
A14.11=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 c5 7.Bb2
A14.12=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 c5 7.Bb2 Nc6
A14.13=Engelskt: Avb�jd Neo-Katalansk, 5...O-O 6.b3 c5 7.Bb2 Nc6 8.e3
A15.1=Engelskt: Engelsk-Indisk
A15.2=Engelskt: Engelsk-Indisk, Polsk
A15.3=Engelskt: Engelsk-Indisk, 2.g3
A15.4=Engelskt: Engelsk-Indisk, 2.g3 e6
A15.5=Engelskt: Engelsk-Indisk, 2.g3 e6 3.Bg2
A15.6=Engelskt: Engelsk-Indisk, 2.g3 g6
A15.7=Engelskt: Engelsk-Indisk, 2.g3 g6 3.Bg2 Bg7
A15.8=Engelskt: Engelsk-Indisk, 2.Nf3
A15.9=Engelskt: Engelsk-Indisk, 2.Nf3 g6
A15.10=Engelskt: Engelsk-Indisk, 2.Nf3 g6 3.g3 Bg7 4.Bg2
A15.11=Engelskt: Engelsk-Indisk, 2.Nf3 g6 3.g3 Bg7 4.Bg2 O-O
A16.1=Engelskt: Engelsk-Indisk, 2.Nc3
A16.2=Engelskt: Engelsk-Indisk, 2.Nc3 Nc6
A16.3=Engelskt: Engelsk-Indisk, 2.Nc3 c6
A16.4=Engelskt: Engelsk-Indisk, 2.Nc3 c6 3.e4
A16.5=Engelskt: Engelsk-Indisk, 2.Nc3 c6 3.e4 d5
A16.7=Engelskt: Engelsk-Indisk, 2.Nc3 d6
A16.8=Engelskt: Engelsk-Indisk, 2.Nc3 g6
A16.9=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.e4
A16.10=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3
A16.11=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7
A16.12=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2
A16.13=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2 O-O
A16.14=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2 O-O 5.e4
A16.15=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2 O-O 5.Nf3
A16.16=Engelskt: Engelsk-Indisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2 O-O 5.Nf3 d6 6.O-O
A16.17=Engelskt: Engelsk-Gr�nfeld
A16.18=Engelskt: Engelsk-Gr�nfeld, 3.Nf3
A16.19=Engelskt: Engelsk-Gr�nfeld, 3.Nf3 g6
A16.20=Engelskt: Engelsk-Gr�nfeld, 3.Nf3 g6 4.Qa4+
A16.21=Engelskt: Engelsk-Gr�nfeld, 3.Nf3 g6 4.g3
A16.22=Engelskt: Engelsk-Gr�nfeld, 3.cxd5
A16.23=Engelskt: Engelsk-Gr�nfeld, Smyslovvarianten
A16.24=Engelskt: Engelsk-Gr�nfeld, Smyslovvarianten, 6.bxc3
A16.25=Engelskt: Engelsk-Gr�nfeld, Smyslovvarianten, 6.bxc3 Bg7
A16.26=Engelskt: Engelsk-Gr�nfeld, Smyslov, 7.Rb1
A16.27=Engelskt: Engelsk-Gr�nfeld, Tjeckisiska varianten
A16.28=Engelskt: Engelsk-Gr�nfeld, 4.Nf3
A16.29=Engelskt: Engelsk-Gr�nfeld, 4.Nf3 g6
A16.30=Engelskt: Engelsk-Gr�nfeld, 4.Nf3 g6 5.g3
A16.31=Engelskt: Engelsk-Gr�nfeld, 4.Nf3 g6 5.g3 Bg7
A16.32=Engelskt: Engelsk-Gr�nfeld, Korchnoivarianten
A16.33=Engelskt: Engelsk-Gr�nfeld, Andersson-B��kvarianten
A16.34=Engelskt: Engelsk-Gr�nfeld, Andersson-B��k, Dambyte
A16.35=Engelskt: Engelsk-Gr�nfeld, 4.Nf3 g6 5.Qa4+
A17.1=Engelskt: Engelsk-Indisk, 2.Nc3 e6
A17.2=Engelskt: Engelsk-Indisk, 2.Nc3 e6 3.g3
A17.3=Engelskt: Engelsk-Indisk, 2.Nc3 e6 3.Nf3
A17.4=Engelskt: Engelsk-Indisk, 2.Nc3 e6 3.Nf3 d5
A17.5=Engelskt: Engelsk-Damindisk
A17.6=Engelskt: Engelsk-Damindisk, 4.e4
A17.7=Engelskt: Engelsk-Damindisk, Romanishin
A17.8=Engelskt: Engelsk-Damindisk, 4.g3
A17.9=Engelskt: Engelsk-Damindisk, 4.g3 Bb7 5.Bg2
A17.10=Engelskt: Engelsk-Damindisk, 4.g3 Bb7 5.Bg2 Be7 6.O-O O-O
A17.11=Engelskt: Engelsk-Damindisk, 4.g3 Bb7 5.Bg2 Be7 6.O-O O-O 7.Re1
A17.12=Engelskt: Nimzo-Engelskt
A17.13=Engelskt: Nimzo-Engelskt, 4.g3
A17.14=Engelskt: Nimzo-Engelskt, 4.Qc2
A17.15=Engelskt: Nimzo-Engelskt, 4.Qc2 O-O
A18.1=Engelskt: Mikenas
A18.2=Engelskt: Mikenas, Kevitz f�rsvar
A18.3=Engelskt: Mikenas, 3...d6
A18.4=Engelskt: Mikenas, Franska varianten
A18.5=Engelskt: Mikenas, Fransk, 4.cxd5
A18.6=Engelskt: Mikenas, Flohrvarianten
A18.7=Engelskt: Mikenas, Flohr, 4...Ne4
A18.8=Engelskt: Mikenas, Flohr, 4...d4
A18.9=Engelskt: Mikenas, Flohr, 7.Nf3
A18.10=Engelskt: Mikenas, Flohr, 7.d4
A19.1=Engelskt: Mikenas, Sicilianska varianten
A19.2=Engelskt: Mikenas, Sicilianskt, 4.e5
A19.3=Engelskt: Mikenas, Sicilianskt, 4.e5 Ng8
A19.4=Engelskt: Mikenas, Neis gambit
A19.5=Engelskt: Mikenas, 5.Nf3
A19.6=Engelskt: Mikenas, 5.Nf3 Nc6
A19.7=Engelskt: Mikenas, 5.Nf3 Nc6 6.d4
A19.8=Engelskt: Mikenas, 6.d4 cxd4 7.Nxd4 Nxe5
A20.1=Engelskt: Avb�jd Kungsindisk, 1...e5
A20.2=Engelskt: Avb�jd Kungsindisk, 2.d3
A20.4=Engelskt: Avb�jd Kungsindisk, 2.g3
A20.5=Engelskt: Avb�jd Kungsindisk, 2.g3 f5
A20.6=Engelskt: Avb�jd Kungsindisk, 2.g3 g6
A20.7=Engelskt: Avb�jd Kungsindisk, 2.g3 g6 3.Bg2
A20.8=Engelskt: Avb�jd Kungsindisk, 2.g3 g6 3.Bg2 Bg7
A20.9=Engelskt: Avb�jd Kungsindisk, 2.g3 c6
A20.10=Engelskt: Avb�jd Kungsindisk, 2.g3 c6 3.d4
A20.11=Engelskt: Avb�jd Kungsindisk, 2.g3 d6
A20.12=Engelskt: Avb�jd Kungsindisk, 2.g3 d6 3.Bg2
A20.13=Engelskt: Avb�jd Kungsindisk, 2.g3 Nc6
A20.14=Engelskt: Avb�jd Kungsindisk, 2.g3 Nc6 3.Bg2
A20.15=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6
A20.16=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6 3.Bg2
A20.17=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6 3.Bg2 Bc5
A20.18=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6 3.Bg2 Nc6
A20.19=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6 3.Bg2 c6
A20.20=Engelskt: Avb�jd Kungsindisk, 2.g3 Nf6 3.Bg2 d5
A20.21=Engelskt: Avb�jd Kungsindisk, Nimzowitsch
A20.22=Engelskt: Avb�jd Kungsindisk, Nimzowitsch, 2...Nc6
A20.23=Engelskt: Avb�jd Kungsindisk, Nimzowitsch, Flohrvarianten
A21.1=Engelskt: Avb�jd Kungsindisk, 2.Nc3
A21.2=Engelskt: Avb�jd Kungsindisk, 2.Nc3 f5
A21.3=Engelskt: Avb�jd Kungsindisk, 2.Nc3 f5 3.g3 Nf6
A21.4=Engelskt: Avb�jd Kungsindisk, 2.Nc3 f5 3.g3 Nf6 4.Bg2
A21.5=Engelskt: Avb�jd Kungsindisk, 2.Nc3 g6
A21.6=Engelskt: Avb�jd Kungsindisk, 2.Nc3 g6 3.g3 Bg7 4.Bg2
A21.7=Engelskt: Avb�jd Kungsindisk, 2.Nc3 d6
A21.8=Engelskt: Avb�jd Kungsindisk, Keresvarianten
A21.9=Engelskt: Avb�jd Kungsindisk, Keresvarianten, 4.Bg2
A21.10=Engelskt: Avb�jd Kungsindisk, 2.Nc3 d6 3.d4
A21.11=Engelskt: Avb�jd Kungsindisk, 2.Nc3 d6 3.g3
A21.12=Engelskt: Avb�jd Kungsindisk, 2.Nc3 d6 3.Nf3
A21.13=Engelskt: Avb�jd Kungsindisk, 2.Nc3 d6 3.Nf3 g6
A21.14=Engelskt: Lukinvarianten
A21.15=Engelskt: Lukin, 4.d4 e4
A21.16=Engelskt: Lukin, 5.Nd2
A21.17=Engelskt: Lukin, 5.Nd2 Nf6 6.e3
A21.18=Engelskt: Lukin, 5.Ng5
A21.19=Engelskt: Lukin, 5.Ng5 Nf6
A21.20=Engelskt: Lukin, 5.Ng5 Be7
A21.21=Engelskt: Lukin, 5.Ng5 c6
A21.22=Engelskt: Smyslovs f�rsvar
A21.23=Engelskt: Kramnik-Shirov motattack
A21.24=Engelskt: Kramnik-Shirov, 3.g3
A21.25=Engelskt: Kramnik-Shirov, 3.g3 Bxc3
A21.26=Engelskt: Kramnik-Shirov, 3.g3 Bxc3 4.bxc3
A21.27=Engelskt: Kramnik-Shirov, 3.Nd5
A21.28=Engelskt: Kramnik-Shirov, 3.Nd5 a5
A21.29=Engelskt: Kramnik-Shirov, 3.Nd5 Ba5
A21.30=Engelskt: Kramnik-Shirov, 3.Nd5 Bc5
A21.31=Engelskt: Kramnik-Shirov, 3.Nd5 Be7
A21.32=Engelskt: Kramnik-Shirov, 3.Nd5 Be7 4.d4
A22.1=Engelskt: Kings, 2.Nc3 Nf6
A22.2=Engelskt: Kings, 2.Nc3 Nf6 3.e4
A22.3=Engelskt: Kings, 2.Nc3 Nf6 3.e3
A22.4=Engelskt: Kings, 2.Nc3 Nf6 3.e3 Bb4
A22.5=Engelskt: Kings, 2.Nc3 Nf6 3.Nf3
A22.6=Engelskt: Kings, 2.Nc3 Nf6 3.Nf3 d6
A22.7=Engelskt: Kings, 2.Nc3 Nf6 3.Nf3 e4
A22.8=Engelskt: Bellons gambit
A22.9=Engelskt: Bremensystemet
A22.10=Engelskt: Bremen, 3...Bc5
A22.11=Engelskt: Bremen, Omv�nd drake
A22.12=Engelskt: Bremen, Omv�nd drake, 4.cxd5
A22.13=Engelskt: Bremen, Omv�nd drake, 4.cxd5 Nxd5
A22.14=Engelskt: Bremen, Omv�nd drake, 4.cxd5 Nxd5 5.Bg2
A22.15=Engelskt: Bremen, Omv�nd drake, 4.cxd5 Nxd5 5.Bg2 Nb6
A22.16=Engelskt: Bremen, Smyslovsystem
A22.17=Engelskt: Bremen, Smyslov, 4.Bg2
A22.18=Engelskt: Bremen, Smyslov, 4.Bg2 Bxc3
A22.19=Engelskt: Bremen, Smyslov, 4.Bg2 O-O
A22.20=Engelskt: Bremen, Smyslov, 4.Bg2 O-O 5.e4
A23.1=Engelskt: Bremen, Keressystem
A23.2=Engelskt: Bremen, Keres, 4.Nf3
A23.3=Engelskt: Bremen, Keres, 4.Nf3 d6
A23.4=Engelskt: Bremen, Keres, 4.Nf3 d6
A23.5=Engelskt: Bremen, Keres, 4.Nf3 e4
A23.6=Engelskt: Bremen, Keres, 4.Bg2
A23.7=Engelskt: Bremen, Keres, 4.Bg2 d5
A23.8=Engelskt: Bremen, Keres, 4.Bg2 d5 5.cxd5
A23.9=Engelskt: Bremen, Keres, 4.Bg2 d5 5.cxd5 cxd5
A24.1=Engelskt: Bremen, 3...g6
A24.2=Engelskt: Bremen, 3...g6 4.Bg2
A24.3=Engelskt: Bremen, 3...g6 4.Bg2 Bg7
A24.4=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.d3
A24.5=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e3
A24.6=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e3 d6 6.Nge2 O-O
A24.7=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e4
A24.8=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e4 d6
A24.9=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e4 d6 6.Nf3
A24.10=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e4 d6 6.Nge2 O-O
A24.11=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.e4 d6 6.Nge2 O-O 7.d3
A24.12=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.Nf3
A24.13=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.Nf3 d6 6.O-O O-O
A24.14=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.Nf3 d6 6.d3 O-O 7.O-O
A24.15=Engelskt: Bremen, 3...g6 4.Bg2 Bg7 5.Nf3 d6 6.d3 O-O 7.O-O c6
A25.1=Engelskt: St�ngd
A25.2=Engelskt: St�ngd, 3.e3
A25.3=Engelskt: St�ngd, 3.e3 Nf6
A25.4=Engelskt: St�ngd, 3.g3
A25.5=Engelskt: St�ngd, 3.g3 f5
A25.6=Engelskt: St�ngd, 3.g3 f5 4.Bg2
A25.7=Engelskt: St�ngd, 3.g3 f5 4.Bg2 Nf6
A25.8=Engelskt: St�ngd, 3.g3 f5 4.Bg2 Nf6 5.e3 g6
A25.9=Engelskt: St�ngd, 3.g3 f5 4.Bg2 Nf6 5.d3
A25.10=Engelskt: St�ngd, 3.g3 Nf6
A25.11=Engelskt: St�ngd, 3.g3 Nf6 4.Bg2
A25.12=Engelskt: St�ngd, 3.g3 Nf6 4.Bg2 Bc5
A25.13=Engelskt: St�ngd, 3.g3 Nf6 4.Bg2 Bc5 5.e3
A25.14=Engelskt: St�ngd, 3.g3 Nf6 4.Bg2 Bb4
A25.15=Engelskt: St�ngd, 3.g3 Nf6 4.Bg2 Bb4 5.Nd5
A25.16=Engelskt: St�ngd, 3.g3 d6 4.Bg2
A25.17=Engelskt: St�ngd, Tr�gers f�rsvar
A25.18=Engelskt: St�ngd, Tr�gers f�rsvar, 5.d3
A25.19=Engelskt: St�ngd, 3.g3 g6
A25.20=Engelskt: St�ngd, 3.g3 g6 4.Bg2
A25.21=Engelskt: St�ngd, 3.g3 g6 4.Bg2 Bg7
A25.22=Engelskt: St�ngd, 3.g6 g6 4.Bg2 Bg7 5.e3
A25.23=Engelskt: St�ngd, Taimanovvarianten
A25.24=Engelskt: St�ngd, Hortvarianten
A25.25=Engelskt: St�ngd, Hortvarianten, 7.d3
A25.26=Engelskt: St�ngd, 5.Rb1
A25.27=Engelskt: St�ngd, 5.Rb1, Taimanovvarianten
A25.28=Engelskt: St�ngd, 5.Rb1 a5
A25.29=Engelskt: St�ngd, 5.e4
A25.30=Engelskt: St�ngd, 5.d3
A25.31=Engelskt: St�ngd, 5.d3 Nge7
A26.1=Engelskt: St�ngd, 5.d3 d6
A26.2=Engelskt: St�ngd, 5.d3 d6 6.e3
A26.3=Engelskt: St�ngd, 5.d3 d6 6.Rb1
A26.4=Engelskt: St�ngd, 5.d3 d6 6.Rb1 f5
A26.5=Engelskt: St�ngd, 5.d3 d6 6.Rb1 a5
A26.6=Engelskt: St�ngd, 5.d3 d6 6.Nf3
A26.7=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6
A26.8=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O
A26.9=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O O-O
A26.10=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O O-O 8.Rb1
A26.11=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O O-O 8.Rb1 a5
A26.12=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O O-O 8.Rb1 a5 9.a3
A26.13=Engelskt: St�ngd, 5.d3 d6 6.Nf3 Nf6 7.O-O O-O 8.Rb1 a5 9.a3 h6
A26.14=Engelskt: Botvinniksystem
A26.15=Engelskt: Botvinniksystem, 6...Nf6
A26.16=Engelskt: Botvinniksystem, 6...Nf6 7.Nf3
A26.17=Engelskt: Botvinniksystem, 6...Nf6 7.Nf3 O-O 8.O-O
A26.18=Engelskt: Botvinniksystem, 6...Nf6 7.Nge2
A26.19=Engelskt: Botvinniksystem, 6...Nf6 7.Nge2 O-O 8.O-O
A26.20=Engelskt: Botvinniksystem, 6...Nge7
A26.21=Engelskt: Botvinniksystem, 6...Nge7 7.Nge2
A27.1=Engelskt: Trespringar
A27.2=Engelskt: Trespringar, 3...Bb4
A27.3=Engelskt: Trespringar, 3...d6
A27.4=Engelskt: Trespringar, 3...f5
A27.5=Engelskt: Trespringar, 3...f5 4.d4
A27.6=Engelskt: Trespringar, 3...f5 4.d4 e4
A27.7=Engelskt: Trespringar, 3...g6
A27.8=Engelskt: Trespringar, 3...g6 4.d4
A27.9=Engelskt: Trespringar, 3...g6 4.d4 exd4
A27.10=Engelskt: Trespringar, 3...g6 4.d4 exd4 5.Nxd4
A28.1=Engelskt: Fyra Springare
A28.2=Engelskt: Fyra Springare, Nimzowitschvarianten
A28.3=Engelskt: Fyra Springare, Marinivarianten
A28.4=Engelskt: Fyra Springare, Capablancavarianten
A28.5=Engelskt: Fyra Springare, 4.d4
A28.6=Engelskt: Fyra Springare, Nenarokovvarianten
A28.7=Engelskt: Fyra Springare, Bradley Beachvarianten
A28.8=Engelskt: Fyra Springare, 4.e3
A28.9=Engelskt: Fyra Springare, 4.e3 Bb4
A28.10=Engelskt: Fyra Springare, 4.e3 Bb4 5.Qc2
A28.11=Engelskt: Fyra Springare, Steanvarianten
A28.12=Engelskt: Fyra Springare, Romanishinvarianten
A29.1=Engelskt: Fyra Springare, 4.g3
A29.2=Engelskt: Fyra Springare, 4.g3 g6
A29.3=Engelskt: Fyra Springare, 4.g3 g6 5.d4
A29.4=Engelskt: Fyra Springare, 4.g3 d5
A29.5=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5
A29.6=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5
A29.7=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2
A29.8=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Be6
A29.9=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6
A29.10=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O
A29.11=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O Be7
A29.12=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O Be7 8.Rb1
A29.13=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O Be7 8.a3
A29.14=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O Be7 8.d3
A29.15=Engelskt: Fyra Springare, 4.g3 d5 5.cxd5 Nxd5 6.Bg2 Nb6 7.O-O Be7 8.d3 O-O
A29.16=Engelskt: Fyra Springare, 4.g3 Bc5
A29.17=Engelskt: Fyra Springare, 4.g3 Bc5 5.Bg2
A29.18=Engelskt: Fyra Springare, 4.g3 Bc5 5.Bg2 d6 6.O-O
A29.19=Engelskt: Fyra Springare, 4.g3 Bc5 5.Bg2 d6 6.O-O O-O
A29.20=Engelskt: Fyra Springare, 4.g3 Bc5 5.Bg2 d6 6.O-O O-O 7.d3
A29.21=Engelskt: Fyra Springare, 4.g3 Bb4
A29.22=Engelskt: Fyra Springare, 4.g3 Bb4 5.Nd5
A29.23=Engelskt: Fyra Springare, 4.g3 Bb4 5.Bg2
A29.24=Engelskt: Fyra Springare, Huvudvarianten 6.O-O
A29.25=Engelskt: Fyra Springare, Huvudvarianten 6.O-O e4
A30.1=Engelskt: Symmetrisk
A30.2=Engelskt: Symmetrisk, 2.b3
A30.3=Engelskt: Symmetrisk, 2.g3
A30.4=Engelskt: Symmetrisk, 2.g3 g6
A30.5=Engelskt: Symmetrisk, 2.Nf3
A30.6=Engelskt: Symmetrisk, 2.Nf3 b6
A30.7=Engelskt: Symmetrisk, 2.Nf3 b6 3.g3
A30.8=Engelskt: Symmetrisk, 2.Nf3 b6 3.g3 Bb7 4.Bg2
A30.9=Engelskt: Symmetrisk, 2.Nf3 g6
A30.10=Engelskt: Symmetrisk, 2.Nf3 Nc6
A30.11=Engelskt: Symmetrisk, 2.Nf3 Nf6
A30.12=Engelskt: Symmetrisk, 2.Nf3 Nf6 3.g3
A30.13=Engelskt: Symmetrisk, b6 System
A30.14=Engelskt: Symmetrisk, b6 System
A30.15=Engelskt: Symmetrisk, b6 System
A30.16=Engelskt: Symmetrisk, b6 system
A30.17=Engelskt: Symmetrisk, Dubbel fianchetto
A30.18=Engelskt: Symmetrisk, Dubbel fianchetto
A30.19=Engelskt: Symmetrisk, �msesidig Dubbelt fianchetto
A30.20=Engelskt: Symmetrisk, �msesidig Dubbelt fianchetto
A30.21=Engelskt: Symmetrisk, �msesidig Dubbelt fianchetto
A30.22=Engelskt: Symmetrisk, �msesidigt Dubbelt fianchetto med ...d5
A30.23=Engelskt: Symmetrisk, Igelkottssystem
A30.24=Engelskt: Symmetrisk, Igelkottssystem
A30.25=Engelskt: Symmetrisk, Igelkottssystem, 6...a6
A30.26=Engelskt: Symmetrisk, Igelkottssystem, 6...d6
A30.27=Engelskt: Symmetrisk, Igelkottssystem, 6...d6 7.b3
A30.28=Engelskt: Symmetrisk, Igelkottssystem, 6...d6 7.d4
A30.29=Engelskt: Symmetrisk, Igelkottssystem
A30.30=Engelskt: Symmetrisk, Igelkottssystem, 7.Re1
A30.31=Engelskt: Symmetrisk, Igelkottssystem, 7.Re1 d5
A30.32=Engelskt: Symmetrisk, Igelkottssystem, 7.b3
A30.33=Engelskt: Symmetrisk, Igelkottssystem, 7.b3
A30.34=Engelskt: Symmetrisk, Igelkottssystem, 7.b3
A30.35=Engelskt: Symmetrisk, Igelkottssystem, 7.d4
A30.36=Engelskt: Symmetrisk, Igelkottssystem, 8.Qxd4
A30.37=Engelskt: Symmetrisk, Igelkottssystem, 8.Qxd4 O-O
A30.38=Engelskt: Symmetrisk, Igelkottssystem, 8.Qxd4 O-O
A30.39=Engelskt: Symmetrisk, Igelkottssystem, 8.Qxd4 Nc6
A30.40=Engelskt: Symmetrisk, Igelkottssystem, 8.Qxd4 d6
A30.41=Engelskt: Symmetrisk, Igelkottssystem, 9.b3
A30.42=Engelskt: Symmetrisk, Igelkottssystem, 9.b3 Nbd7
A30.43=Engelskt: Symmetrisk, Igelkottssystem, 9.b3 Nbd7 10.Nb5
A30.44=Engelskt: Symmetrisk, Igelkottssystem, 9.Rd1
A30.45=Engelskt: Symmetrisk, Igelkottssystem, Flexibel formation
A30.46=Engelskt: Symmetrisk, Igelkottssystem, Flexibel formation
A30.47=Engelskt: Symmetrisk, Igelkottssystem, Flexibel formation, 11.e4 Qc7
A30.48=Engelskt: Symmetrisk, Igelkottssystem, Flexibel formation, 11.e4 O-O
A31.1=Engelskt: Symmetrisk, Tv� springare, 1.c4 c5 2.Nf3 Nf6 3.d4
A31.2=Engelskt: Symmetrisk, Tv� springare, 3...a6
A31.3=Engelskt: Symmetrisk, Tv� springare, 3...g6
A31.4=Engelskt: Symmetrisk, Tv� springare, 3...g6 4.d5
A31.5=Engelskt: Symmetrisk, Tv� springare, 3...g6 4.Nc3
A31.6=Engelskt: Symmetrisk, Tv� springare, 3..cxd4
A31.7=Engelskt: Symmetrisk, Tv� springare, 3..cxd4 4.Nxd4
A31.8=Engelskt: Symmetrisk, Tv� springare, 4...b6
A31.9=Engelskt: Symmetrisk, Tv� springare, 4...b6 5.Nc3 Bb7
A31.10=Engelskt: Symmetrisk, Tv� springare, 4...g6
A31.11=Engelskt: Symmetrisk, Tv� springare, 4...g6 5.Nc3
A31.12=Engelskt: Symmetrisk, Tv� springare, 4...g6 5.Nc3 Bg7
A31.13=Engelskt: Symmetrisk, Tv� springare, 4...g6
A31.14=Engelskt: Symmetrisk, Tv� springare, 4...Nc6
A31.15=Engelskt: Symmetrisk, Tv� springare, 4...Nc6 5.Nc3
A31.16=Engelskt: Symmetrisk, Tv� springare, 4...Nc6 5.Nc3 g6
A31.17=Engelskt: Symmetrisk, Tv� springare, 4...e5
A31.18=Engelskt: Symmetrisk, Tv� springare, 4...e5 5.Nb5
A32.1=Engelskt: Symmetrisk, Tv� springare, 4...e6
A32.2=Engelskt: Symmetrisk, Tv� springare, 5.e3
A32.3=Engelskt: Symmetrisk, Tv� springare, 5.g3
A32.4=Engelskt: Symmetrisk, Tv� springare, 5.g3 a6
A32.5=Engelskt: Symmetrisk, Tv� springare, 5.g3 a6
A32.6=Engelskt: Symmetrisk, Tv� springare, 5.g3 Qb6
A32.7=Engelskt: Symmetrisk, Tv� springare, 5.g3 Qb6 6.Bg2
A32.8=Engelskt: Symmetrisk, Tv� springare, 5.g3 Qc7
A32.9=Engelskt: Symmetrisk, Tv� springare, 5.g3 Nc6
A32.10=Engelskt: Symmetrisk, Tv� springare, 5.g3 Nc6 6.Bg2
A32.11=Engelskt: Symmetrisk, Tv� springare, 5.g3 Bb4+
A32.12=Engelskt: Symmetrisk, Tv� springare, 5.g3 d5
A32.15=Engelskt: Symmetrisk, Tv� springare, 5.Nc3
A32.16=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 d5
A32.17=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 a6
A32.18=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 a6 6.g3
A32.19=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Bb4
A32.20=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Bb4 6.Qb3
A32.21=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Bb4 6.Nb5
A32.22=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Bb4 6.Bd2
A32.23=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Bb4 6.Bd2 Nc6
A33.1=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6
A33.2=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Bf4
A33.3=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Bg5
A33.4=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.e3
A33.5=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.a3
A33.6=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.a3 Bc5
A33.7=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Ndb5
A33.8=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Ndb5 Bb4
A33.9=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Ndb5 d5
A33.10=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.Ndb5 d5 Dambyte
A33.11=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.g3
A33.12=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.g3 a6
A33.13=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.g3 Bb4
A33.14=Engelskt: Symmetrisk, Tv� springare, 5.Nc3 Nc6 6.g3 Bc5
A33.15=Engelskt: Symmetrisk, Gellervarianten
A33.16=Engelskt: Symmetrisk, Geller, 7.Nb3
A33.17=Engelskt: Symmetrisk, Geller, 7.Nb3 Ne5
A34.1=Engelskt: Symmetrisk
A34.2=Engelskt: Symmetrisk, 2...b6
A34.3=Engelskt: Symmetrisk, 2...b6 3.Nf3
A34.4=Engelskt: Symmetrisk, 2...b6 3.Nf3 Bb7
A34.5=Engelskt: Symmetrisk, 2...g6
A34.6=Engelskt: Symmetrisk, 2...g6 3.Nf3
A34.7=Engelskt: Symmetrisk, 2...g6 3.g3
A34.8=Engelskt: Symmetrisk, 2...g6 3.g3 Bg7 4.Bg2
A34.9=Engelskt: Symmetrisk, 2...Nf6
A34.11=Engelskt: Symmetrisk, 2...Nf6 3.g3
A34.10=Engelskt: Symmetrisk, 2...Nf6 3.g3 d5
A34.12=Engelskt: Symmetrisk, 2...Nf6 3.g3 d5 4.cxd5 Nxd5 5.Bg2
A34.13=Engelskt: Symmetrisk, Rubinsteinsystemet
A34.14=Engelskt: Symmetrisk, Tre springare
A34.15=Engelskt: Symmetrisk, Tre springare, 3...b6
A34.16=Engelskt: Symmetrisk, Tre springare, 3...e6
A34.17=Engelskt: Symmetrisk, Tre springare, 3...e6 4.g3
A34.18=Engelskt: Symmetrisk, Tre springare, 3...g6
A34.19=Engelskt: Symmetrisk, Tre springare
A34.20=Engelskt: Symmetrisk, Tre springare, Avbyte
A34.21=Engelskt: Symmetrisk, Tre springare, 5.g3
A34.22=Engelskt: Symmetrisk, Tre springare, 5.e4
A34.23=Engelskt: Symmetrisk, Tre springare, 5.e4 Nxc3
A34.24=Engelskt: Symmetrisk, Tre springare, Dambyte
A34.25=Engelskt: Symmetrisk, Tre springare, 5.e4 Nb4
A34.26=Engelskt: Symmetrisk, Tre springare, 5.e4 Nb4 6.Bb5+
A34.27=Engelskt: Symmetrisk, Tre springare, 5.e4 Nb4 6.Bc4
A34.28=Engelskt: Symmetrisk, Tre springare, 5.d4
A34.29=Engelskt: Symmetrisk, Tre springare, 5.d4 cxd4
A34.30=Engelskt: Symmetrisk, Tre springare, 5.d4 Nxc3
A35.1=Engelskt: Symmetrisk
A35.2=Engelskt: Symmetrisk, 2.Nc3 Nc6 3.e3
A35.3=Engelskt: Symmetrisk, 2.Nc3 Nc6 3.Nf3
A35.4=Engelskt: Symmetrisk, 2.Nc3 Nc6 3.Nf3 g6
A35.5=Engelskt: Symmetrisk, 2.Nc3 Nc6 3.Nf3 g6 4.e3
A35.6=Engelskt: Symmetrisk, 2.Nc3 Nc6 3.Nf3 g6 4.e3 Bg7
A35.7=Engelskt: Symmetrisk, Fyra Springare
A35.8=Engelskt: Symmetrisk, Fyra Springare, 4.d4
A35.9=Engelskt: Symmetrisk, Fyra Springare, 4.e3
A35.10=Engelskt: Symmetrisk, Fyra Springare, 4.e3 e5
A35.11=Engelskt: Symmetrisk, Fyra Springare, 4.g3
A35.12=Engelskt: Symmetrisk, Fyra Springare, 4.g3 d5
A35.13=Engelskt: Symmetrisk, Fyra Springare, 4.g3 d5 5.cxd5
A36.1=Engelskt: Symmetrisk, 3.g3
A36.2=Engelskt: Symmetrisk, 3.g3 Nf6
A36.3=Engelskt: Symmetrisk, 3.g3 e6
A36.4=Engelskt: Symmetrisk, 3.g3 e6 4.Nf3
A36.5=Engelskt: Symmetrisk, Keres-Parmasystemet
A36.6=Engelskt: Symmetrisk, Keres-Parma, Huvudvarianten Avbyte
A36.7=Engelskt: Symmetrisk, 3.g3 g6
A36.8=Engelskt: Symmetrisk, 3.g3 g6 4.Bg2
A36.9=Engelskt: Symmetrisk, 3.g3 g6 4.Bg2 Bg7
A36.10=Engelskt: Symmetrisk, 5.d3
A36.11=Engelskt: Symmetrisk, 5.a3
A36.12=Engelskt: Symmetrisk, 5.a3 e6
A36.13=Engelskt: Symmetrisk, 5.a3 d6
A36.14=Engelskt: Symmetrisk, 5.b3
A36.15=Engelskt: Symmetrisk, 5.e3
A36.16=Engelskt: Symmetrisk, 5.e3 e5 (Botvinnik Omv�nd)
A36.17=Engelskt: Symmetrisk, 5.e3 e6
A36.18=Engelskt: Symmetrisk, 5.e3 e6 6.Nge2
A36.19=Engelskt: Symmetrisk, 5.e3 e6 6.Nge2 Nge7
A36.20=Engelskt: Symmetriskt, Botvinniksystem
A36.21=Engelskt: Symmetriskt, Botvinniksystem, 5...Nf6
A36.22=Engelskt: Symmetriskt, Botvinniksystem, 5...Nf6 6.Nge2
A36.23=Engelskt: Symmetriskt, Botvinniksystem, 5...e6
A36.24=Engelskt: Symmetriskt, Botvinniksystem, 5...e6 6.Nge2 Nge7
A36.25=Engelskt: Symmetriskt, Botvinniksystem, 5...e6, 8.d3
A36.26=Engelskt: Symmetriskt, Botvinniksystem, 5...e6, 8.d3 d6
A36.27=Engelskt: Symmetriskt, Botvinniksystem, 5...d6
A36.28=Engelskt: Symmetriskt, Botvinniksystem, 5...d6 6.Nge2
A36.29=Engelskt: Symmetriskt, Botvinniksystem, 5...d6 6.Nge2 Nf6
A36.30=Engelskt: Symmetriskt, Botvinniksystem, 5...d6, 7.O-O O-O
A36.31=Engelskt: Symmetriskt, Botvinniksystem, 5...d6, 8.d3
A36.32=Engelskt: Symmetriskt, Botvinniksystem, 5...d6, 8.d3 Rb8
A36.33=Engelskt: Symmetriskt, Botvinniksystem, 5...d6, 8.d3 Ne8
A36.34=Engelskt: Symmetriskt, Botvinniksystem, 5...d6, 8.d3 a6
A37.1=Engelskt: Symmetrisk, 5.Nf3
A37.2=Engelskt: Symmetrisk, 5.Nf3 a6
A37.3=Engelskt: Symmetrisk, 5.Nf3 Nh6
A37.4=Engelskt: Symmetrisk, 5.Nf3 Nh6 6.O-O
A37.5=Engelskt: Symmetrisk, 5.Nf3 d6
A37.6=Engelskt: Symmetrisk, 5.Nf3 d6 6.d3
A37.7=Engelskt: Symmetrisk, 5.Nf3 d6 6.O-O
A37.8=Engelskt: Symmetrisk, 5.Nf3 d6 6.O-O Nh6
A37.9=Engelskt: Symmetrisk, 5.Nf3 e6
A37.10=Engelskt: Symmetrisk, 5.Nf3 e6 6.d3
A37.11=Engelskt: Symmetrisk, 5.Nf3 e6 6.e3
A37.12=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O
A37.13=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O Nge7
A37.14=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O Nge7 7.e3
A37.15=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O Nge7 7.d3
A37.16=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O Nge7 7.d3 O-O
A37.17=Engelskt: Symmetrisk, 5.Nf3 e6 6.O-O Nge7 7.d3 O-O 8.Bd2
A37.18=Engelskt: Symmetrisk, 5.Nf3 e5
A37.19=Engelskt: Symmetrisk, 5.Nf3 e5 6.a3
A37.20=Engelskt: Symmetrisk, 5.Nf3 e5 6.d3
A37.21=Engelskt: Symmetrisk, 5.Nf3 e5 6.d3 Nge7
A37.22=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O
A37.23=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O d6
A37.24=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O d6 7.d3
A37.25=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O d6 7.d3 Nge7
A37.26=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O d6 7.d3 Nge7 8.a3
A37.27=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O Nge7
A37.28=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O Nge7 7.d3
A37.29=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O Nge7 7.d3 O-O
A37.30=Engelskt: Symmetrisk, 5.Nf3 e5 6.O-O Nge7 7.d3 O-O 8.a3
A38.1=Engelskt: Symmetrisk, Huvudvarianten
A38.2=Engelskt: Symmetrisk, Huvudvarianten, 6.d4
A38.3=Engelskt: Symmetrisk, Huvudvarianten, 6.O-O
A38.4=Engelskt: Symmetrisk, Huvudvarianten, 6.O-O d5
A38.5=Engelskt: Symmetrisk, Huvudvarianten, 6.O-O d6
A38.6=Engelskt: Symmetrisk, Huvudvarianten, 6.O-O O-O
A38.7=Engelskt: Symmetrisk, Huvudvarianten, 7.Rb1
A38.8=Engelskt: Symmetrisk, Huvudvarianten, 7.b3
A38.9=Engelskt: Symmetrisk, Huvudvarianten, 7.a3
A38.10=Engelskt: Symmetrisk, Huvudvarianten, 7.a3 d6
A38.11=Engelskt: Symmetrisk, Huvudvarianten, 7.d3
A38.12=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 a6
A38.13=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d5
A38.14=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d6
A38.15=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d6 8.Rb1
A38.16=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d6 8.Bd2
A38.17=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d6 8.a3
A38.18=Engelskt: Symmetrisk, Huvudvarianten, 7.d3 d6 8.a3 a6
A39.1=Engelskt: Symmetrisk, Huvudvarianten 7.d4
A39.2=Engelskt: Symmetrisk, Huvudvarianten 7.d4 cxd4
A39.3=Engelskt: Symmetrisk, Huvudvarianten 7.d4 cxd4 8.Nxd4
A39.4=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Qa5
A39.5=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Qb6
A39.6=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Qb6
A39.7=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...a6
A39.8=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...d6
A39.9=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Ng4
A39.10=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Ng4 9.e3 d6
A39.11=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 8...Nxd4
A39.12=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 9.Qxd4
A39.13=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 9...d6
A39.14=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd2
A39.15=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3
A39.16=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 Bf5
A39.17=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 Rb8
A39.18=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 a6
A39.19=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 a6 11.Bd2
A39.20=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 a6 11.Bd2 Rb8
A39.21=Engelskt: Symmetrisk, Huvudvarianten 7.d4, 10.Qd3 a6 11.Bd2 Rb8 12.Rac1
A40.1=Dambondeparti
A40.2=Dambonde: 1...c6
A40.3=Dambonde: 1...c6 2.Nf3
A40.4=Dambonde: 1...c6 2.c4
A40.5=Dambonde: Jadoul
A40.6=Dambonde: Polskt f�rsvar
A40.7=Dambonde: Polskt f�rsvar
A40.8=Dambonde: Polskt f�rsvar
A40.9=Dambonde: Polskt f�rsvar, Spasskys gambit
A40.10=Dambonde: Engelskt f�rsvar
A40.11=Dambonde: Engelskt f�rsvar, 2.c4
A40.12=Dambonde: Engelskt f�rsvar, 2.c4 Bb7
A40.13=Dambonde: Engelskt f�rsvar, 2.c4 e6
A40.14=Dambonde: Engelskt f�rsvar, 3.a3
A40.15=Dambonde: Engelskt f�rsvar, 3.e4
A40.16=Dambonde: Engelskt f�rsvar, Pollis gambit
A40.17=Dambonde: Engelskt f�rsvar, Hartlaubs gambit
A40.18=Dambonde: Engelskt f�rsvar, 3.Nc3
A40.19=Englunds (Charlick) gambit
A40.20=Antagen Englunds (Charlick) gambit
A40.21=Englunds (Charlick) gambit: Soller
A40.22=Englunds (Charlick) gambit: Hartlaub
A40.23=Englunds (Charlick) gambit: 2.dxe5 Nc6
A40.24=Englunds (Charlick) gambit: 2.dxe5 Nc6 3.Nf3
A40.25=Englunds (Charlick) gambit: Avb�jd Soller
A40.26=Englunds (Charlick) gambit: Zilbermints
A40.27=Englunds (Charlick) gambit: 2.dxe5 Nc6 3.Nf3 Qe7
A40.28=Dambonde: Lundins (Kevitz-Mikenas-Bogoljubow-Miles) f�rsvar
A40.29=Dambonde: Bogoljubow-Miles, 2.Bg5
A40.30=Dambonde: Bogoljubow-Miles, 2.d5
A40.31=Dambonde: Bogoljubow-Miles, 2.c4
A40.32=Dambonde: Bogoljubow-Miles, Pozareks gambit
A40.33=Dambonde: Bogoljubow-Miles, 2.Nf3
A40.34=Dambonde: 1...e6
A40.35=Dambonde: 1...e6 2.Nf3
A40.37=Dambonde: 1...e6 2.c4
A40.38=Dambonde: Keres f�rsvar
A40.39=Dambonde: Keres f�rsvar, 3.Bd2
A40.40=Dambonde: Keres f�rsvar, 3.Bd2 Bxd2+
A40.41=Dambonde: Keres f�rsvar, K�ngru-varianten
A40.42=Dambonde: Keres f�rsvar, 3.Bd2 a5
A40.43=Dambonde: Modern, 1.d4 g6
A40.44=Dambonde: Modern, 1.d4 g6 2.Nf3
A40.45=Dambonde: Modern, 1.d4 g6 2.c4
A40.46=Dambonde: Modern, 1.d4 g6 2.c4 Bg7
A40.47=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.e4
A40.48=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.Nf3
A40.49=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.Nf3 c5
A40.50=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.Nc3
A40.51=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.Nc3 c5
A40.52=Dambonde: Modern, 1.d4 g6 2.c4 Bg7 3.Nc3 c5 4.d5
A40.53=Dambonde: Modern, Beefeaters f�rsvar
A41.1=Neo-Gammalindisk
A41.2=Neo-Gammalindiskt: 2.Bg5
A41.3=Neo-Gammalindiskt: 2.g3
A41.4=Neo-Gammalindiskt: 2.Nf3
A41.5=Neo-Gammalindiskt: Modern
A41.6=Neo-Gammalindiskt: Modern, 3.Bf4
A41.7=Neo-Gammalindiskt: Modern, 3.Bf4 Bg7
A41.8=Neo-Gammalindiskt: Modern, 3.g3
A41.9=Neo-Gammalindiskt: Modern, 3.g3 Bg7
A41.10=Neo-Gammalindiskt: Modern, 3.g3 Bg7 4.Bg2
A41.11=Neo-Gammalindiskt: Wades f�rsvar
A41.12=Neo-Gammalindiskt: Wades f�rsvar, 3.e3
A41.13=Neo-Gammalindiskt: Wades f�rsvar, 3.e3 Nd7
A41.14=Neo-Gammalindiskt: Wades f�rsvar, 3.e3 Nf6
A41.15=Neo-Gammalindiskt: Wades f�rsvar, 3.c4
A41.16=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 e5
A41.17=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 e5 4.Nc3
A41.18=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 e5 4.Nc3 Nc6
A41.19=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 e5 4.dxe5
A41.20=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 e5 4.dxe5 Nc6 gambit
A41.21=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 Nd7
A41.22=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 Nd7 4.Nc3
A41.24=Neo-Gammalindiskt: Wades f�rsvar, 3.c4 Bxf3
A41.25=Neo-Gammalindiskt: Wades f�rsvar, 3.e4
A41.26=Neo-Gammalindiskt: Wades f�rsvar, 3.e4 Nf6
A41.27=Neo-Gammalindiskt: 2.c4
A41.28=Neo-Gammalindiskt: 2.c4 e5
A41.29=Neo-Gammalindiskt: 2.c4 e5 3.d5
A41.30=Neo-Gammalindiskt: 2.c4 e5 3.dxe5
A41.31=Neo-Gammalindiskt: Dambyte
A41.32=Neo-Gammalindiskt: 2.c4 e5 3.Nf3
A41.33=Neo-Gammalindiskt: 2.c4 e5 3.Nf3 e4
A41.34=Neo-Gammalindiskt: Modern, 2.c4 g6
A41.35=Neo-Gammalindiskt: Modern, 3.e4
A41.36=Neo-Gammalindiskt: Modern, 3.e4 Bg7
A41.37=Neo-Gammalindiskt: Modern, 3.Nf3
A41.38=Neo-Gammalindiskt: Modern, 3.Nf3 Bg7
A41.39=Neo-Gammalindiskt: Modern, 3.Nf3 Bg7 4.g3
A41.40=Neo-Gammalindiskt: Modern, 3.Nf3 Bg7 4.e4
A41.41=Neo-Gammalindiskt: Modern, Rossolimovarianten
A41.42=Neo-Gammalindiskt: Modern, 3.Nc3
A41.43=Neo-Gammalindiskt: Modern, 3.Nc3 Bg7
A41.44=Neo-Gammalindiskt: Modern, 3.Nc3 Bg7 4.Nf3
A41.45=Neo-Gammalindiskt: Modern, 3.Nc3 Bg7 4.Nf3 Bf4
A41.46=Neo-Gammalindiskt: Modern, 3.Nc3 Bg7 4.Nf3 Bf4 5.e3
A41.47=Neo-Gammalindiskt: Modern, 3.Nc3 Bg7 4.Nf3 Bf4 5.e3 Nc6
A42.1=Moderna: Averbakh
A42.2=Moderna: Averbakh, Randspringervarianten
A42.3=Moderna: Averbakh, Randspringer, 5.Nf3
A42.4=Moderna: c4 Pterodactyl
A42.5=Moderna: c4 Pterodactyl, 5.Nf3
A42.6=Moderna: c4 Pterodactyl, 5.Nf3 Qa5
A42.7=Moderna: Averbakh, 4...c6
A42.8=Moderna: Averbakh, 4...c6 5.Be3
A42.9=Moderna: Averbakh, 4...c6 5.Nf3
A42.10=Moderna: Averbakh, 4...Nd7
A42.11=Moderna: Averbakh, 4...Nd7 5.Nf3
A42.12=Moderna: Averbakh, Kotovvarianten
A42.13=Moderna: Averbakh, Kotov, 5.Nf3
A42.14=Moderna: Averbakh, Kotov, 5.Nge2
A42.15=Moderna: Averbakh, Kotov, 5.d5
A42.16=Moderna: Averbakh, Kotov, 5.Be3
A42.17=Moderna: Averbakh, Kotov, 5.Be3 e5
A42.18=Moderna: Averbakh, Kotov, 5.Be3 e5 6.Nge2
A42.19=Moderna: Averbakh, Kotov, 5.Be3 e5 6.d5
A42.20=Moderna: Averbakh, Kotov, 5.Be3 e5 6.d5 Nce7
A42.21=Moderna: Averbakh, Kotov, 5.Be3 e5 6.d5 Nce7 7.c5
A42.22=Moderna: Averbakh, Kotov, 5.Be3 e5 6.d5 Nce7 7.g4
A42.23=Moderna: Averbakh, 4...e5
A42.24=Moderna: Averbakh, 4...e5 5.Nge2
A42.25=Moderna: Averbakh, 4...e5 5.Nf3
A42.26=Moderna: Averbakh, 4...e5 5.Nf3 Nd7
A42.27=Moderna: Averbakh, 4...e5 5.Nf3 Nd7 6.Be2
A42.28=Moderna: Averbakh, 4...e5 5.Nf3 Nd7 6.Be2 Ne7
A42.29=Moderna: Averbakh, 4...e5 5.d5
A42.30=Moderna: Averbakh, 4...e5 5.d5 Nd7
A42.31=Moderna: Averbakh, 4...e5 5.dxe5
A42.32=Moderna: Averbakh, 4...e5 5.dxe5 dxe5
A42.33=Moderna: Averbakh, Dambyte
A42.34=Moderna: Averbakh, Dambyte, 7.f4
A43.1=Gamla Benoni
A43.2=Gamla Benoni: Nakamuras gambit
A43.3=Gamla Benoni: 2.dxc5
A43.4=Gamla Benoni: Cormorants gambit
A43.5=Gamla Benoni: 2.c3
A43.6=Gamla Benoni: 2.e3
A43.7=Gamla Benoni: 2.d5
A43.8=Gamla Benoni: 2.d5 b5
A43.9=Gamla Benoni: 2.d5 e6
A43.10=Gamla Benoni: Franco-Benoni
A43.11=Gamla Benoni: 2.d5 e6 3.c4
A43.12=Gamla Benoni: 2.d5 e6 3.c4
A43.13=Gamla Benoni: 2.d5 e6 3.c4
A43.14=Gamla Benoni: 2.d5 e6 3.c4
A43.15=Gamla Benoni: 2.d5 e6 3.c4
A43.16=Gamla Benoni: 2.d5 e6 3.c4
A43.17=Gamla Benoni: 2.d5 e6 3.c4
A43.18=Gamla Benoni: Clarendon Court f�rsvar
A43.19=Gamla Benoni: 2.d5 Nf6
A43.20=Gamla Benoni: 2.d5 Nf6 3.Nc3
A43.21=Gamla Benoni: Woozle
A43.22=Gamla Benoni: 2.d5 Nf6 3.Nf3
A43.23=Gamla Benoni: 2.d5 Nf6 3.Nf3 e6
A43.24=Gamla Benoni: 2.d5 Nf6 3.Nf3 e6 4.Nc3
A43.25=Gamla Benoni: 2.d5 Nf6 3.Nf3 g6
A43.26=Gamla Benoni: 2.d5 Nf6 3.Nf3 g6 4.Nc3
A43.27=Gamla Benoni: Neo-Benko
A43.28=Gamla Benoni: Neo-Benko, 4.Bg5
A43.29=Gamla Benoni: Neo-Benko, 4.Bg5 d6
A43.30=Gamla Benoni: Neo-Benko, 4.Bg5 Ne4
A43.31=Gamla Benoni: Hawk
A43.32=Gamla Benoni: Hawk, 4.e4
A43.33=Gamla Benoni: Schmidt
A43.34=Gamla Benoni: Schmidt, 3.Nf3
A43.35=Gamla Benoni: Schmidt, 3.Nf3 Nf6
A43.36=Gamla Benoni: Schmidt, 3.Nc3
A43.37=Gamla Benoni: Schmidt, 3.Nc3 g6
A43.38=Gamla Benoni: Schmidt, 3.Nc3 Nf6
A43.39=Gamla Benoni: Schmidt, 3.e4
A43.40=Gamla Benoni: Schmidt, 3.e4 g6
A43.41=Gamla Benoni: Schmidt, 3.e4 g6
A43.42=Gamla Benoni: Schmidt, 3.e4 g6
A43.43=Gamla Benoni: Schmidt, 3.e4 g6
A43.44=Gamla Benoni: Schmidt, 3.e4 Nf6
A43.45=Gamla Benoni: Schmidt, 3.e4 Nf6
A43.46=Gamla Benoni: Schmidt, 3.e4 Nf6
A43.47=Gamla Benoni: Schmidt, 3.e4 Nf6
A43.48=Gamla Benoni: Schmidt, 3.e4 Nf6
A43.49=Gamla Benoni: Schmidt, 6.h3
A43.50=Gamla Benoni: Schmidt, 6.h3
A43.51=Gamla Benoni: Schmidt, 6.Bb5+
A43.52=Gamla Benoni: Schmidt, 6.Be2
A43.53=Gamla Benoni: Schmidt, 6.Be2 O-O
A43.54=Gamla Benoni: Schmidt, 6.Be2 O-O 7.O-O
A43.55=Gamla Benoni: Schmidt, 6.Be2 O-O 7.O-O e6
A43.56=Gamla Benoni: Schmidt, 6.Be2 O-O 7.O-O Na6
A43.57=Gamla Benoni: Schmidt, 6.Be2 O-O 7.O-O Na6 8.h3
A44.1=Gamla Benoni: Tjeckiskt
A44.2=Gamla Benoni: Tjeckiskt, 3.dxe6
A44.3=Gamla Benoni: Tjeckiskt, 3.c4
A44.4=Gamla Benoni: Tjeckiskt, 3.c4 d6
A44.5=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4
A44.6=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 Be7
A44.7=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 Be7 5.Nc3
A44.8=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 g6
A44.9=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 g6 5.Nc3
A44.10=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 g6 5.Nc3 Bg7
A44.11=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 g6 5.Nc3 Bg7 6.Nf3
A44.12=Gamla Benoni: Tjeckiskt, 3.c4 d6 4.e4 g6 5.Nc3 Bg7 6.Bd3
A44.13=Gamla Benoni: Tjeckiskt, 3.e4
A44.14=Gamla Benoni: Tjeckiskt, 3.e4 d6
A44.15=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nf3
A44.16=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Bb5+
A44.17=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Bd3
A44.18=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3
A44.19=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 Nf6
A44.20=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 g6
A44.21=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 a6
A44.22=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 a6 5.a4 Be7
A44.23=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 Be7
A44.24=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 Be7 5.Bb5+
A44.25=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 Be7 5.Nf3
A44.26=Gamla Benoni: Tjeckiskt, 3.e4 d6 4.Nc3 Be7 5.Nf3 Bg4
A45.1=Dambonde: Indian
A45.2=Indiskt: Blekansikte-attack
A45.3=Indiskt: Blackmar-Diemers gambit (utan Nc3)
A45.4=Indiskt: T�lamodsattack
A45.5=Indiskt: Omegas gambit
A45.6=Indiskt: Arafats gambit
A45.7=Indiskt: Gibbins gambit
A45.8=Indiskt: Gibbins gambit, Oshima f�rsvar
A45.9=Indiskt: Antagen Gibbins gambit
A45.10=Indiskt: Canard �ppning
A45.11=Indiskt: 2.Nd2
A45.12=Indiskt: Lazards gambit
A45.13=Indiskt: 2.e3
A45.14=Indiskt: 2.e3 e6
A45.15=Indiskt: 2.e3 g6
A45.16=Indiskt: 2.c3
A45.17=Indiskt: 2.c3 g6
A45.18=Indiskt: 2.c3 g6 3.Bg5
A45.19=Indiskt: 2.Nc3
A45.20=Indiskt: 2.Bf4
A45.21=Indiskt: 2.g3
A45.22=Indiskt: 2.g3 g6
A45.23=Indiskt: 2.g3 c5
A45.24=Indiskt: 2.g3 c5 3.d5 b5
A45.25=Trompowskys �ppning
A45.26=Trompowsky 2...d6
A45.27=Trompowsky 2...d6 3.Nc3
A45.28=Trompowsky 2...d6 3.Bxf6
A45.29=Trompowsky 2...g6
A45.30=Trompowsky 2...g6 3.Nc3
A45.31=Trompowsky 2...g6 3.Bxf6
A45.32=Trompowsky 2...g6 3.Bxf6 exf6 4.e3
A45.33=Trompowsky: 2...e6
A45.34=Trompowsky: 2...e6 3.Nc3
A45.35=Trompowsky: 2...e6 3.e3
A45.36=Trompowsky: 2...e6 3.Nd2
A45.37=Trompowsky: 2...e6 3.e4
A45.38=Trompowsky: 2...e6 3.e4 h6
A45.39=Trompowsky: 2...e6 3.e4 h6 4.Bxf6
A45.40=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6
A45.41=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.c3
A45.42=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.Nc3
A45.43=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.Nc3 Bb4
A45.44=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.Nc3 d6
A45.45=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.Nc3 d6 6.Qd2
A45.46=Trompowsky: 2...e6 3.e4 h6 4.Bxf6 Qxf6 5.Nc3 d6 6.Qd2 g5
A45.47=Trompowsky: 2...c5
A45.48=Trompowsky: 2...c5 3.dxc5
A45.49=Trompowsky: 2...c5 3.Nc3
A45.50=Trompowsky: 2...c5 3.d5
A45.51=Trompowsky: 2...c5 3.d5 Qb6
A45.52=Trompowsky: 2...c5 3.d5 Qb6 4.Nc3
A45.53=Trompowsky: 2...c5 3.Bxf6
A45.54=Trompowsky: 2...c5 3.Bxf6 gxf6
A45.55=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5
A45.56=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6
A45.57=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1
A45.58=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1 f5
A45.59=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1 f5 6.c4
A45.60=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1 f5 6.g3
A45.61=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1 f5 6.e3
A45.62=Trompowsky: 2...c5 3.Bxf6 gxf6 4.d5 Qb6 5.Qc1 f5 6.e3 Bg7
A45.63=Trompowsky: 2...Ne4
A45.64=Trompowsky: 2...Ne4 3.h4
A45.65=Trompowsky: 2...Ne4 3.h4 d5
A45.66=Trompowsky: 2...Ne4 3.h4 c5
A45.67=Trompowsky: 2...Ne4 3.h4 c5 4.dxc5
A45.68=Trompowsky: 2...Ne4 3.h4 c5 4.d5
A45.69=Trompowsky: 2...Ne4 3.Bh4
A45.70=Trompowsky: 2...Ne4 3.Bh4 g5
A45.71=Trompowsky: 2...Ne4 3.Bh4 d5
A45.72=Trompowsky: 2...Ne4 3.Bh4 c5
A45.73=Trompowsky: 2...Ne4 3.Bh4 c5 4.f3
A45.74=Trompowsky: 2...Ne4 3.Bf4
A45.75=Trompowsky: Borgvarianten
A45.76=Trompowsky: 2...Ne4 3.Bf4 d5
A45.77=Trompowsky: 2...Ne4 3.Bf4 d5 4.Nd2
A45.78=Trompowsky: 2...Ne4 3.Bf4 d5 4.f3
A45.79=Trompowsky: 2...Ne4 3.Bf4 d5 4.f3 Nf6
A45.80=Trompowsky: 2...Ne4 3.Bf4 d5 4.e3
A45.81=Trompowsky: 2...Ne4 3.Bf4 d5 4.e3 c5
A45.82=Trompowsky: 2...Ne4 3.Bf4 c5
A45.83=Trompowsky: 2...Ne4 3.Bf4 c5 4.d5
A45.84=Trompowsky: 2...Ne4 3.Bf4 c5 4.d5 Qb6
A45.85=Trompowsky: 2...Ne4 3.Bf4 c5 4.f3
A45.86=Trompowsky: 2...Ne4 3.Bf4 c5 4.f3 Qa5+
A45.87=Trompowsky: 2...Ne4 3.Bf4 c5 4.f3 Qa5+ 5.c3 Nf6 6.d5
A45.88=Trompowsky: 2...Ne4 3.Bf4 c5 4.f3 Qa5+ 5.c3 Nf6 6.Nd2
A46.1=Indiskt: 2.Nf3
A46.2=Indiskt: D�rys f�rsvar
A46.3=Indiskt: 2.Nf3 b5
A46.4=Indiskt: 2.Nf3 b5 3.g3
A46.5=Neo-Benoni
A46.6=Neo-Benoni 3.dxc5
A46.7=Neo-Benoni: 3.e3
A46.8=Neo-Benoni: 3.e3 cxd4
A46.9=Neo-Benoni: 3.c3
A46.10=Neo-Benoni: 3.c3 cxd4
A46.11=Neo-Benoni: 3.c3 b6
A46.12=Neo-Benoni: 3.c3 g6
A46.13=Neo-Benoni: 3.c3 e6
A46.14=Neo-Benoni: 3.g3
A46.15=Neo-Benoni: 3.g3 cxd4
A46.16=Neo-Benoni: 3.g3 cxd4 4.Nxd4
A46.17=Indiskt: 2.Nf3 d6
A46.18=Indiskt: 2.Nf3 d6 3.g3
A46.19=Indiskt: 2.Nf3 d6 3.Bg5
A46.20=Indiskt: 2.Nf3 d6 3.Bg5 Nbd7
A46.21=Indiskt: 2.Nf3 e6
A46.22=Indiskt: 2.Nf3 e6 3.c3
A46.23=Indiskt: 2.Nf3 e6 3.c3 b6
A46.24=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.c3 b6 4.Bg5
A46.25=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.e3
A46.26=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.e3 c5
A46.27=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.e3 c5 4.Bd3
A46.28=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3
A46.29=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 b5
A46.30=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 b5 4.Bg2 Bb7
A46.31=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 b5 4.Bg2 Bb7 5.O-O
A46.32=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5
A46.33=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5 4.Bg2
A46.34=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5 4.Bg2 cxd4
A46.35=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5 4.Bg2 Nc6
A46.36=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5 4.Bg2 Qc7
A46.37=Indiskt: 1.d4 Nf6 2.Nf3 e6 3.g3 c5 4.Bg2 Qa5+
A46.38=Indiskt: Londonsystem
A46.39=Indiskt: London, 3...c5
A46.40=Indiskt: London, 3...c5 4.e3
A46.41=Indiskt: London, 3...c5 4.e3 Qb6
A46.42=Indiskt: London, 3...c5 4.c3
A46.43=Torreattack
A46.44=Torreattack: 3...b6
A46.45=Torreattack: 3...Be7
A46.46=Torreattack: 3...c5
A46.47=Torreattack: Wagners gambit
A46.48=Torreattack: 3...c5 4.c3
A46.49=Torreattack: 3...c5 4.c3 Qb6
A46.50=Torreattack: 3...c5 4.c3 h6
A46.51=Torreattack: 3...c5 4.c3 h6 5.Bh4
A46.52=Torreattack: 3...c5 4.e3
A46.53=Torreattack: 3...c5 4.e3 cxd4
A46.54=Torreattack: 3...c5 4.e3 Qb6
A46.55=Torreattack: 3...c5 4.e3 Be7
A46.56=Torreattack: 3...c5 4.e3 h6
A46.57=Torreattack: 3...c5 4.e3 h6 5.Bh4
A46.58=Torreattack: 3...h6
A46.59=Torreattack: 3...h6 4.Bh4
A46.60=Torreattack: 3...h6 4.Bh4 g5
A46.61=Torreattack: 3...h6 4.Bxf6
A46.62=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4
A46.63=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 b6
A46.64=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 c5
A46.65=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 d6
A46.66=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 d6 6.Nc3
A46.67=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 d6 6.Nc3 g6
A46.68=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 d6 6.Nc3 Nd7
A46.69=Torreattack: 3...h6 4.Bxf6 Qxf6 5.e4 d6 6.Nc3 Nd7 7.Qd2
A47.1=Neo-Damindiskt 1.d4 Nf6 2.Nf3 b6
A47.2=Neo-Damindiskt 2..b6 3.Bf4
A47.3=Neo-Damindiskt 2..b6 3.Bf4 e6
A47.4=Neo-Damindiskt 2..b6 3.Bf4 e6 4.e3
A47.5=Neo-Damindiskt 2..b6 3.Bf4 e6 4.e3 c5
A47.6=Neo-Damindiskt 2..b6 3.Bf4 Bb7
A47.7=Neo-Damindiskt 2..b6 3.Bf4 Bb7 4.e3
A47.8=Neo-Damindiskt 2..b6 3.Bf4 Bb7 4.e3 e6
A47.9=Neo-Damindiskt 2..b6 3.Bg5
A47.10=Neo-Damindiskt 2..b6 3.Bg5 Bb7
A47.11=Neo-Damindiskt 2..b6 3.e3
A47.12=Neo-Damindiskt 2..b6 3.e3 e6
A47.13=Neo-Damindiskt 2..b6 3.e3 e6 4.Bd3
A47.14=Neo-Damindiskt 2..b6 3.e3 e6 4.Bd3 c5
A47.15=Neo-Damindiskt 2..b6 3.e3 Bb7
A47.16=Neo-Damindiskt 2..b6 3.e3 Bb7 4.Bd3
A47.17=Neo-Damindiskt 2..b6 3.e3 Bb7 4.Bd3 e6
A47.18=Neo-Damindiskt 2..b6 3.e3 Bb7 4.Bd3 e6 5.O-O
A47.19=Neo-Damindiskt 2..b6 3.e3 Bb7 4.Bd3 e6 5.O-O c5
A47.20=Neo-Damindiskt 2..b6 3.g3
A47.21=Neo-Damindiskt 2..b6 3.g3 e6
A47.22=Neo-Damindiskt 2..b6 3.g3 Bb7 4.Bg2
A47.23=Neo-Damindiskt 2..b6 3.g3 Bb7 4.Bg2 e6
A47.24=Neo-Damindiskt Marienbadsystemet
A47.25=Neo-Damindiskt Marienbadsystemet, Bergvarianten
A48.1=Neo-Kungsindiskt: �stindiskt f�rsvar, 1.d4 Nf6 2.Nf3 g6
A48.2=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.Nbd2
A48.3=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.c3
A48.4=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.c3 Bg7
A48.5=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.e3
A48.6=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.e3 Bg7
A48.7=Neo-Kungsindiskt: �stindiskt f�rsvar, 2..g6 3.e3 c5
A48.8=Neo-Kungsindiskt: �stindiskt f�rsvar, 1.d4 Nf6 2.Nf3 g6 3.Nc3
A48.9=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4
A48.10=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7
A48.11=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.Nbd2
A48.12=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.c3
A48.13=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.e3
A48.14=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.e3 O-O
A48.15=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.e3 O-O 5.Be2
A48.16=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.e3 O-O 5.Be2 d6
A48.17=Neo-Kungsindiskt: Londonsystemet,  2..g6 3.Bf4 Bg7 4.e3 O-O 5.Be2 d6 6.h3
A48.18=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5
A48.19=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Ne4
A48.20=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7
A48.21=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.c3
A48.22=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.e3
A48.23=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nc3
A48.24=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2
A48.25=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O
A48.26=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.e4
A48.27=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.e4 d6
A48.28=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.e4 d5
A48.29=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.c3
A48.30=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.c3 d6
A48.31=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.c3 d6 6.e4
A48.32=Neo-Kungsindiskt: Torreattack,  2..g6 3.Bg5 Bg7 4.Nbd2 O-O 5.c3 d6 6.e4 c5
A49.1=Neo-Kungsindiskt: Fianchettosystemet, 1.d4 Nf6 2.Nf3 g6 3.g3
A49.2=Neo-Kungsindiskt: Fianchettosystemet, 2..g6 3.g3 Bg7
A49.3=Neo-Kungsindiskt: Fianchettosystemet, 2..g6 3.g3 Bg7 4.Bg2
A49.4=Neo-Kungsindiskt: Fianchettosystemet, 2..g6 3.g3 Bg7 4.Bg2 O-O
A49.5=Neo-Kungsindiskt: Dubbla Fianchettosystemet, 2..g6 3.g3 Bg7 4.Bg2 O-O 5.b3 d6 6.Bb2
A49.6=Neo-Kungsindiskt: Fianchettosystemet, 2..g6 3.g3 Bg7 4.Bg2 O-O 5.O-O
A49.7=Neo-Kungsindiskt: Fianchettosystemet, 2..g6 3.g3 Bg7 4.Bg2 O-O 5.O-O d6
A50.1=Indiskt: 2.c4
A50.2=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar)
A50.3=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nc3
A50.4=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nf3
A50.5=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nf3 d6
A50.6=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nf3 e6
A50.7=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nf3 e6 4.a3
A50.8=Indiskt: Svart springartango (Mexikanskt f�rsvar-Kevitz-Trajkovich f�rsvar), 3.Nf3 e6 4.Nc3
A50.9=Indiskt: Slavisk-Indisk, 1.d4 Nf6 2.c4 c6
A50.10=Indiskt: Slavisk-Indisk, 1.d4 Nf6 2.c4 c6 3.Nf3 3.Nf3
A50.11=Indiskt: Slavisk-Indisk, 1.d4 Nf6 2.c4 c6 3.Nc3 3.Nc3
A50.12=Indiskt: 2.c4 a6
A50.13=Indiskt: Damindisk Accelererad, 1.d4 Nf6 2.c4 b6
A50.14=Indiskt: Damindisk Accelererad, 1.d4 Nf6 2.c4 b6 3.Nc3 Bb7
A50.15=Indiskt: Damindisk Accelererad, 1.d4 Nf6 2.c4 b6 3.Nc3 Bb7 4.Qc2
A51.1=Budapestf�rsvaret
A51.2=Budapestf�rsvaret: 3.e3
A51.3=Budapestf�rsvaret: 3.d5
A51.4=Budapestf�rsvaret: 3.dxe5
A51.5=Budapestf�rsvaret: Fajarowicz-Richters gambit
A51.6=Budapestf�rsvaret: Fajarowicz-Richters gambit, Steinervarianten
A51.7=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.Nd2
A51.8=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.a3
A51.9=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.Nf3
A51.10=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.Nf3 Bb4+
A51.11=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.Nf3 Nc6
A51.12=Budapestf�rsvaret: Fajarowicz-Richters gambit, 4.Nf3 Nc6 5.a3
A52.1=Budapestf�rsvaret: 3...Ng4
A52.2=Budapestf�rsvaret: 3...Ng4 4.e3
A52.3=Budapestf�rsvaret: Alekhinevarianten
A52.4=Budapestf�rsvaret: Alekhinevarianten, Baloghs gambit
A52.5=Budapestf�rsvaret: Alekhinevarianten, Abonyivarianten
A52.6=Budapestf�rsvaret: Adlervarianten
A52.7=Budapestf�rsvaret: Adler, 4...Bc5
A52.8=Budapestf�rsvaret: Adler, 4...Bc5 5.e3 Nc6 6.Be2
A52.9=Budapestf�rsvaret: Rubinsteinvarianten
A52.10=Budapestf�rsvaret: Rubinstein, 4...Bb4+
A52.11=Budapestf�rsvaret: Rubinstein, 4...Nc6
A52.12=Budapestf�rsvaret: Rubinstein, Huvudvarianten
A52.13=Budapestf�rsvaret: Rubinstein, Huvudvarianten, 6.Nbd2
A52.14=Budapestf�rsvaret: Rubinstein, Huvudvarianten, 6.Nbd2 Qe7 7.e3
A53.1=Gammalindiskt
A53.2=Gammalindiskt: 3.g3
A53.3=Gammalindiskt: 3.Nf3
A53.4=Gammalindiskt: 3.Nf3 c6
A53.5=Gammalindiskt: 3.Nf3 Nbd7
A53.6=Gammalindiskt: 3.Nf3 Bf5
A53.7=Gammalindiskt: 3.Nf3 Bg4
A53.8=Gammalindiskt: 3.Nf3 Bg4 4.Qb3
A53.9=Gammalindiskt: 3.Nf3 Bg4 4.Nc3
A53.10=Gammalindiskt: 3.Nc3
A53.11=Gammalindiskt: 3.Nc3 c6
A53.12=Gammalindiskt: 3.Nc3 Nbd7
A53.13=Gammalindiskt: 3.Nc3 Nbd7 4.Nf3
A53.14=Gammalindiskt: 3.Nc3 Nbd7 4.e4
A53.15=Gammalindiskt: 3.Nc3 Nbd7 4.e4 e5
A53.16=Gammalindiskt: 3.Nc3 Nbd7 4.e4 e5 5.d5
A53.17=Gammalindiskt: 3.Nc3 Nbd7 4.e4 e5 5.Nge2
A53.18=Gammalindiskt: Janowski
A53.19=Gammalindiskt: Ukrainsk
A53.20=Gammalindiskt: Ukrainsk, 4.e4
A53.21=Gammalindiskt: Ukrainsk, 4.e3
A53.22=Gammalindiskt: Dus-Khotimirsky
A53.23=Gammalindiskt: Ukrainsk, 4.d5
A53.24=Gammalindiskt: Ukrainsk, 4.d5 Be7
A53.25=Gammalindiskt: Ukrainsk, 4.dxe5
A53.26=Gammalindiskt: Ukrainsk, Dambyte
A53.27=Gammalindiskt: Ukrainsk, Dambyte, 6.Nf3
A53.28=Gammalindiskt: Ukrainsk, Dambyte, 6.Nf3 Nfd7
A54.1=Gammalindiskt: 4.Nf3
A54.2=Gammalindiskt: 4.Nf3 exd4
A54.3=Gammalindiskt: 4.Nf3 Nc6
A54.4=Gammalindiskt: 4.Nf3 e4
A54.5=Gammalindiskt: 4.Nf3 e4 5.Ng5
A54.6=Gammalindiskt: 4.Nf3 Nbd7
A54.7=Gammalindiskt: 5.e3
A54.8=Gammalindiskt: 5.g3
A54.9=Gammalindiskt: 5.g3 c6
A54.10=Gammalindiskt: 5.g3 c6 6.Bg2
A54.11=Gammalindiskt: 5.g3 g6
A54.12=Gammalindiskt: 5.g3 g6 6.Bg2
A54.13=Gammalindiskt: 5.g3 g6 6.Bg2 Bg7
A54.14=Gammalindiskt: 5.g3 Be7
A54.15=Gammalindiskt: 5.g3 Be7 6.Bg2
A54.16=Gammalindiskt: 5.g3 Be7 6.Bg2 O-O
A54.17=Gammalindiskt: 5.g3 Be7 6.Bg2 O-O 7.O-O
A54.18=Gammalindiskt: 5.g3 Be7, Huvudvarianten
A54.19=Gammalindiskt: 5.g3 Be7, Huvudvarianten, 8.Qc2
A54.20=Gammalindiskt: 5.Bg5
A54.21=Gammalindiskt: 5.Bg5 c6
A54.22=Gammalindiskt: 5.Bg5 Be7
A54.23=Gammalindiskt: 5.Bg5 Be7 6.e3
A54.24=Gammalindiskt: 5.Bg5 Be7 6.e3 c6
A54.25=Gammalindiskt: 5.Bg5 Be7 6.e3 O-O
A54.26=Gammalindiskt: 5.Bg5 Be7 6.e3 O-O 7.Qc2
A54.27=Gammalindiskt: 5.Bg5 Be7 6.e3 O-O 7.Qc2 c6
A55.1=Gammalindiskt: 5.e4
A55.2=Gammalindiskt: 5.e4 g6
A55.3=Gammalindiskt: 5.e4 c6
A55.4=Gammalindiskt: 5.e4 c6 6.Be2
A55.5=Gammalindiskt: 5.e4 Be7
A55.6=Gammalindiskt: 5.e4 Be7 6.g3
A55.7=Gammalindiskt: 5.e4 Be7 6.g3 O-O
A55.8=Gammalindiskt: 5.e4 Be7 6.g3 c6
A55.9=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2
A55.10=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O
A55.11=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O 8.O-O
A55.12=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O 8.O-O Qc7
A55.13=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O 8.O-O Re8
A55.14=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O 8.O-O a6
A55.15=Gammalindiskt: 5.e4 Be7 6.g3 c6 7.Bg2 O-O 8.O-O a6 9.a4
A55.16=Gammalindiskt: 5.e4 Be7 6.Be2
A55.17=Gammalindiskt: 5.e4 Be7 6.Be2 O-O
A55.18=Gammalindiskt: 5.e4 Be7 6.Be2 c6
A55.19=Gammalindiskt: 5.e4 Be7 6.Be2 c6 7.O-O
A55.20=Gammalindiskt: 5.e4 Be7 6.Be2 c6 7.O-O a6
A55.21=Gammalindiskt: Huvudvarianten
A55.22=Gammalindiskt: Huvudvarianten, 8.h3
A55.23=Gammalindiskt: Huvudvarianten, 8.Be3
A55.24=Gammalindiskt: Huvudvarianten, 8.Be3 a6
A55.25=Gammalindiskt: Huvudvarianten, 8.Qc2
A55.26=Gammalindiskt: Huvudvarianten, 8.Qc2 Re8
A55.27=Gammalindiskt: Huvudvarianten, 8.Qc2 Qc7
A55.28=Gammalindiskt: Huvudvarianten, 8.Qc2 a6
A55.29=Gammalindiskt: Huvudvarianten, 8.Re1
A55.30=Gammalindiskt: Huvudvarianten, 8.Re1 Re8
A55.31=Gammalindiskt: Huvudvarianten, 8.Re1 a6
A55.32=Gammalindiskt: Huvudvarianten, 8.Re1 a6 9.Bf1
A56.1=Benoni: 2...c5
A56.2=Benoni: 2...c5 3.e3
A56.3=Benoni: 2...c5 3.e3 e6
A56.4=Benoni: 2...c5 3.e3 g6
A56.5=Benoni: 2...c5 3.e3 g6 4.Nc3
A56.6=Benoni: 3.dxc5
A56.7=Benoni: 3.d5
A56.8=Benoni: 3.d5 a6
A56.9=Benoni: 3.d5 g6
A56.10=Benoni: 3.d5 g6 4.Nc3
A56.11=Benoni: 3.d5 d6
A56.12=Benoni: 3.d5 d6 4.Nc3 g6
A56.13=Benoni: Bronsteins gambit
A56.14=Benoni: 3.d5 d6 4.Nc3 g6 5.e4 Bg7
A56.17=Benoni: Vulture
A56.18=Benoni: Tjeckiskt
A56.19=Benoni: Tjeckiskt, 4.Nc3 d6
A56.20=Benoni: Tjeckiskt, 5.e4 g6
A56.21=Benoni: Tjeckiskt, 5.e4 Be7
A56.22=Benoni: Tjeckiskt, 5.e4 Be7 6.g3
A56.23=Benoni: Tjeckiskt, 5.e4 Be7 6.g3 O-O
A56.24=Benoni: Tjeckiskt, 5.e4 Be7 6.g3 O-O 7.Bg2
A56.25=Benoni: Tjeckiskt, 5.e4 Be7 6.g3 O-O 7.Bg2 Ne8
A56.26=Benoni: Tjeckiskt, 5.e4 Be7 6.Bd3
A56.27=Benoni: Tjeckiskt, 5.e4 Be7 6.Nf3
A56.28=Benoni: Tjeckiskt, 5.e4 Be7 6.Nf3 O-O
A56.29=Benoni: Tjeckiskt, 5.e4 Be7 6.Nf3 O-O 7.h3
A56.30=Benoni: Tjeckiskt, 5.e4 Be7 6.Nf3 O-O 7.Be2
A57.1=Benkogambit
A57.2=Benkogambit: 4.a4
A57.3=Benkogambit: 4.Nd2
A57.4=Benkogambit: 4.Nf3
A57.5=Benkogambit: 4.Nf3 bxc4
A57.6=Benkogambit: 4.Nf3 Bb7
A57.7=Benkogambit: 4.Nf3 Bb7 5.a4
A57.8=Benkogambit: 4.Nf3 g6
A57.9=Benkogambit: 4.Nf3 g6 5.cxb5
A57.10=Benkogambit: 4.Nf3 g6 5.cxb5 a6
A57.11=Benkogambit: 4.cxb5
A57.12=Benkogambit: 4.cxb5 a6
A57.13=Benkogambit: 4.cxb5 a6 5.b6
A57.14=Benkogambit: 4.cxb5 a6 5.b6 Qxb6
A57.15=Benkogambit: 4.cxb5 a6 5.b6 d6
A57.16=Benkogambit: 4.cxb5 a6 5.b6 e6
A57.17=Benkogambit: 4.cxb5 a6 5.e3
A57.18=Benkogambit: 4.cxb5 a6 5.e3 g6
A57.19=Benkogambit: 4.cxb5 a6 5.e3 g6 6.Nc3 d6
A57.20=Benkogambit: 4.cxb5 a6 5.e3 g6 6.Nc3 Bg7
A57.21=Benkogambit: 4.cxb5 a6 5.f3
A57.22=Benkogambit: 4.cxb5 a6 5.f3 e6
A57.23=Benkogambit: 4.cxb5 a6 5.f3 axb5
A57.24=Benkogambit: Zaitsevvarianten
A57.25=Benkogambit: Zaitsev, 5...Qa5
A57.26=Benkogambit: Zaitsev, 5...axb5
A57.27=Benkogambit: Zaitsev, 5...axb5 6.e4 b4
A57.28=Benkogambit: Zaitsev, 8.Nf3
A57.29=Benkogambit: Zaitsev, Nescafe Frappe attack
A57.30=Benkogambit: Zaitsev, 8.Bf4
A57.31=Benkogambit: Zaitsev, 8.Bf4 g5
A58.1=Benkogambit: 5.bxa6
A58.2=Benkogambit: 5.bxa6 g6
A58.3=Benkogambit: 5.bxa6 Bxa6
A58.4=Benkogambit: Antagen, 6.g3
A58.5=Benkogambit: Antagen, 6.g3 d6 7.Bg2 g6
A58.6=Benkogambit: Antagen, 6.g3 d6 7.Bg2 g6 8.b3
A58.7=Benkogambit: Antagen, 6.Nc3
A58.8=Benkogambit: Antagen, 6.Nc3 g6
A58.9=Benkogambit: Antagen, 6.Nc3 d6
A58.10=Benkogambit: Antagen, 7.f4
A58.11=Benkogambit: Antagen, 7.f4
A58.12=Benkogambit: Antagen, 7.g3
A58.13=Benkogambit: Antagen, 7.g3
A58.14=Benkogambit: Antagen, 7.Nf3
A58.15=Benkogambit: Antagen, 7.Nf3 g6
A58.16=Benkogambit: Antagen, 7.Nf3 g6 8.Nd2
A58.17=Benkogambit: Antagen, 7.Nf3 g6 8.Nd2 Qa5
A58.18=Benkogambit: Antagen, 7.Nf3 g6 8.Nd2 Bg7
A58.19=Benkogambit: Fianchettovarianten, 7.Nf3 g6 8.g3
A58.20=Benkogambit: Fianchettovarianten, 7.Nf3 g6 8.g3 Bg7
A58.21=Benkogambit: Fianchetto, 9.Bh3
A58.22=Benkogambit: Fianchetto, 9.Bg2
A58.23=Benkogambit: Fianchetto, 9...Nbd7
A58.24=Benkogambit: Fianchetto, 9...Nbd7 10.O-O Nb6
A58.25=Benkogambit: Fianchetto, 9...O-O
A58.26=Benkogambit: Fianchetto, Huvudvarianten
A58.27=Benkogambit: Fianchetto, Huvudvarianten, 11.Rb1
A58.28=Benkogambit: Fianchetto, Huvudvarianten, 11.Re1
A58.29=Benkogambit: Fianchetto, Huvudvarianten, 11.Qc2
A58.30=Benkogambit: Fianchetto, Huvudvarianten, 11.Qc2 Qb6
A59.1=Benkogambit: 7.e4
A59.2=Benkogambit: 7.e4 Bxf1 8.Kxf1 g6
A59.3=Benkogambit: 7.e4 Line, 9.Nge2
A59.4=Benkogambit: 7.e4 Line, 9.Nf3
A59.5=Benkogambit: 7.e4 Line, 9.Nf3 Bg7 10.h3
A59.6=Benkogambit: 7.e4 Line, 9.Nf3 Bg7 10.h3 Nbd7
A59.7=Benkogambit: 7.e4 Line, 9.g4
A59.8=Benkogambit: 7.e4 Line, 9.g3
A59.9=Benkogambit: 7.e4, Huvudvarianten
A59.10=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7
A59.11=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.Re1
A59.12=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.Re1 Qa5
A59.13=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.Re1 Ng4
A59.14=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3
A59.15=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Ra6
A59.16=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Ra6 13.Re1
A59.17=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Qb6
A59.18=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Qb6 13.Re1
A59.19=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Qa5
A59.20=Benkogambit: 7.e4, Huvudvarianten, 11...Nbd7 12.h3 Qa5 13.Re1
A60.1=Benoni: 3.d5 e6
A60.2=Benoni: 4.Nf3
A60.3=Benoni: 4.Nf3 exd5 5.cxd5
A60.4=Benoni: Ormvarianten mot 4.Nf3
A60.5=Benoni: 4.g3
A60.6=Benoni: 4.g3 exd5 5.cxd5 b5
A60.7=Benoni: 4.Nc3
A60.8=Benoni: 4.Nc3 exd5 5.Nxd5
A60.9=Benoni: 4.Nc3 exd5 5.cxd5
A60.10=Benoni: Ormvarianten
A60.11=Benoni: Ormen, 6.Nf3
A60.12=Benoni: Ormen, 6.Nf3 Bc7
A60.13=Benoni: Ormen, 6.e4
A60.14=Benoni: Ormen, 6.e4 O-O 7.Nf3
A60.15=Benoni: 4.Nc3 exd5 5.cxd5 g6
A60.16=Benoni: 4.Nc3 exd5 5.cxd5 d6
A60.17=Benoni: 4.Nc3 exd5 5.cxd5 d6 6.Nf3
A61.1=Benoni: 6.Nf3 g6
A61.2=Benoni: 6.Nf3 g6 7.h3
A61.3=Benoni: 6.Nf3 g6 7.Bf4
A61.4=Benoni: 6.Nf3 g6 7.Bf4 a6
A61.5=Benoni: 6.Nf3 g6 7.Bf4 Bg7
A61.6=Benoni: 6.Nf3 g6 7.Bf4 Bg7 8.Nd2
A61.7=Benoni: 6.Nf3 g6 7.Bf4 Bg7 8.Qa4+
A61.8=Benoni: Uhlmannvarianten
A61.9=Benoni: Uhlmann, 7...Bg7
A61.10=Benoni: Uhlmann, 7...h6
A61.11=Benoni: Nimzowitschvarianten
A61.12=Benoni: Nimzowitschvarianten, 7...Nbd7
A61.13=Benoni: Nimzowitschvarianten, 7...Bg7
A61.14=Benoni: Nimzowitschvarianten, 7...Bg7 8.Nc4 O-O 9.Bf4
A61.15=Benoni: Nimzowitschvarianten, 7...Bg7 8.Nc4 O-O 9.Bg5
A61.16=Benoni: Fianchettovarianten
A62.1=Benoni: Fianchettovarianten, 8.Bg2 O-O
A62.2=Benoni: Fianchettovarianten, 9.O-O
A62.3=Benoni: Fianchettovarianten, 9.O-O a6
A62.4=Benoni: Fianchettovarianten, 9.O-O Na6
A62.5=Benoni: Fianchettovarianten, 9.O-O Na6 10.Nd2 Nc7
A62.6=Benoni: Fianchettovarianten, 9.O-O Re8
A63.1=Benoni: Fianchettovarianten, 9...Nbd7
A63.2=Benoni: Fianchettovarianten, 9...Nbd7 10.Nd2
A63.3=Benoni: Fianchettovarianten, 9...Nbd7 10.Nd2 Re8
A63.4=Benoni: Fianchettovarianten, 9...a6 10.a4 Nbd7
A63.5=Benoni: Fianchettovarianten, 9...Nbd7 10.Nd2 a6
A63.6=Benoni: Fianchettovarianten, 9...Nbd7 10.Nd2 a6 11.a4
A64.1=Benoni: Fianchetto, 11...Re8
A64.2=Benoni: Fianchetto, 11...Re8 12.a5
A64.3=Benoni: Fianchetto, 11...Re8 12.Nc4
A64.4=Benoni: Fianchetto, 11...Re8 12.Nc4 Ne5
A64.5=Benoni: Fianchetto, 11...Re8 12.h3
A64.6=Benoni: Fianchetto, 11...Re8 12.h3 Rb8
A64.7=Benoni: Fianchetto, 11...Re8 12.h3 Rb8 13.Nc4
A64.8=Benoni: Fianchetto, 11...Re8 12.h3 Rb8 13.Nc4 Ne5
A64.9=Benoni: Fianchetto, 11...Re8 12.h3 Rb8 13.Nc4 Nb6
A65.1=Benoni: 6.e4
A65.2=Benoni: 6.e4 Be7
A65.3=Benoni: 6.e4 g6
A65.4=Benoni: 6.e4 g6 7.h3
A65.5=Benoni: 6.e4 g6 7.Bf4
A65.8=Benoni: 6.e4 g6 7.Bf4 a6 8.Nf3 b5 9.Qe2
A65.9=Benoni: 6.e4 g6 7.Bd3
A65.10=Benoni: 6.e4 g6 7.Bd3 Bg7 8.h3
A65.11=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2
A65.12=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2 O-O
A65.13=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2 O-O 9.O-O
A65.14=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2 O-O 9.O-O b6
A65.15=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2 O-O 9.O-O Na6
A65.16=Benoni: 6.e4 g6 7.Bd3 Bg7 8.Nge2 O-O 9.O-O a6
A65.17=Benoni: S�misch (6.e4 g6 7.f3)
A65.18=Benoni: S�misch, 7...Bg7
A65.19=Benoni: S�misch, 8.Nge2
A65.20=Benoni: S�misch, 8.Be3
A65.21=Benoni: S�misch, 8.Bg5
A65.22=Benoni: S�misch, 8.Bg5 O-O
A65.23=Benoni: S�misch, 8.Bg5 O-O 9.Nge2
A65.24=Benoni: S�misch, 8.Bg5 O-O 9.Qd2
A65.25=Benoni: S�misch, 8.Bg5 O-O 9.Qd2 a6
A65.26=Benoni: S�misch, 8.Bg5 h6
A65.27=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O
A65.28=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Nge2
A65.29=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2
A65.30=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 Re8
A65.31=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6
A65.32=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6 11.a4
A65.33=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6 11.a4 h5
A65.34=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6 11.a4 Nbd7
A65.35=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6 11.a4 Re8
A65.36=Benoni: S�misch, 8.Bg5 h6 9.Be3 O-O 10.Qd2 a6 11.a4 Re8 12.Nge2 Nbd7
A66.1=Benoni: Fyrbondeattack, 1.d4 Nf6 2.c4 c5 3.d5 e6 4.Nc3 exd5 5.cxd5 d6 6.e4 g6 7.f4
A66.2=Benoni: Fyrbondeattack, 7.f4 Bg7
A66.3=Benoni: Fyra b�nder, Mikenas attack
A66.4=Benoni: Mikenas attack, 8...dxe5
A66.5=Benoni: Mikenas attack, 8...Nfd7
A66.6=Benoni: Mikenas attack, 8...Nfd7 9.e6
A66.7=Benoni: Mikenas attack, 8...Nfd7 9.Nf3
A66.8=Benoni: Mikenas attack, 8...Nfd7 9.Nb5
A66.9=Benoni: Mikenas attack, 9.Nb5 dxe5 10.Nd6+
A66.10=Benoni: Mikenas attack, 9.Nb5 dxe5 10.Nd6+ Ke7 11.Nxc8+
A66.11=Benoni: Mikenas attack, 9.Nb5 dxe5 10.Nd6+ Ke7 11.Nxc8+ Qxc8 12.Nf3
A67.1=Benoni: Fyra b�nder, Taimanov (Alatortsev)varianten
A67.2=Benoni: Fyra b�nder, Taimanov, 8...Nbd7
A67.3=Benoni: Fyra b�nder, Taimanov, 8...Nbd7 9.e5 dxe5 10.fxe5 Nh5 11.e6
A67.4=Benoni: Fyra b�nder, Taimanov, 8...Nfd7
A67.5=Benoni: Fyra b�nder, Taimanov, 9.Bd3
A67.6=Benoni: Fyra b�nder, Taimanov, 9.Bd3 O-O
A67.7=Benoni: Fyra b�nder, Taimanov, 9.Bd3 O-O 10.Nf3
A67.8=Benoni: Fyra b�nder, Taimanov, 9.Bd3 O-O 10.Nf3 a6
A67.9=Benoni: Fyra b�nder, Taimanov, 9.Bd3 O-O 10.Nf3 a6
A67.10=Benoni: Fyra b�nder, Taimanov, 9.Bd3 O-O 10.Nf3 Na6
A67.11=Benoni: Fyra b�nder, Taimanov, 9.a4 (Zaitsev)
A67.12=Benoni: Fyra b�nder, Taimanov, 9.a4 Qh4+
A67.13=Benoni: Fyra b�nder, Taimanov, 9.a4 a6
A67.14=Benoni: Fyra b�nder, Taimanov, 9.a4 a6 10.Bd3
A67.15=Benoni: Fyra b�nder, Taimanov, 9.a4 a6 10.Be2
A67.16=Benoni: Fyra b�nder, Taimanov, 9.a4 O-O
A67.17=Benoni: Fyra b�nder, Taimanov, 9.a4 O-O 10.Nf3
A67.18=Benoni: Fyra b�nder, Taimanov, 9.a4 O-O 10.Nf3 Na6
A67.19=Benoni: Fyra b�nder, Taimanov, 9.a4 O-O 10.Nf3 Na6 11.O-O Nc7
A68.1=Benoni: Fyra b�nder, 8.Nf3
A68.2=Benoni: Fyra b�nder, 8.Nf3 O-O
A68.3=Benoni: Fyra b�nder, 9.Bd3
A68.4=Benoni: Fyra b�nder, 9.Be2
A68.5=Benoni: Fyra b�nder, 9.Be2 b5
A68.6=Benoni: Fyra b�nder, 9.Be2 b5 10.e5
A68.7=Benoni: Fyra b�nder, 9.Be2 b5 10.e5 dxe5
A68.8=Benoni: Fyra b�nder, 9.Be2 b5 10.e5 dxe5 11.fxe5 Ng4 12.Bg5
A68.9=Benoni: Fyra b�nder, 9.Be2 Bg4
A68.10=Benoni: Fyra b�nder, 9.Be2 Bg4 10.e5
A68.11=Benoni: Fyra b�nder, 9.Be2 Bg4 10.O-O
A68.12=Benoni: Fyra b�nder, 9.Be2 Bg4 10.O-O Nbd7
A68.13=Benoni: Fyra b�nder, 9.Be2 Bg4 10.O-O Nbd7 11.h3
A68.14=Benoni: Fyra b�nder, 9.Be2 Bg4 10.O-O Nbd7 11.h3 Bxf3 12.Bxf3 Re8
A68.15=Benoni: Fyra b�nder, 9.Be2 Bg4 10.O-O Nbd7 11.h3 Bxf3 12.Bxf3 Re8 13.Re1
A69.1=Benoni: Fyra b�nder, Huvudvarianten
A69.2=Benoni: Fyra b�nder, Huvudvarianten, 10.O-O
A69.3=Benoni: Fyra b�nder, Huvudvarianten, 10.Nd2
A69.4=Benoni: Fyra b�nder, Huvudvarianten, 10.Nd2 a6
A69.5=Benoni: Fyra b�nder, Huvudvarianten, 10.Nd2 Nbd7
A69.6=Benoni: Fyra b�nder, Huvudvarianten, 10.e5
A69.7=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.O-O
A69.8=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.e6
A69.9=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.Bg5
A69.10=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.Bg5 f6
A69.11=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.Bg5 Qb6
A69.12=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.Bg5 Qb6 13.O-O Nxe5 14.Nxe5
A69.13=Benoni: Fyra b�nder, Huvudvarianten, 10.e5: 12.Bg5 Qb6 13.O-O Nxe5 14.d6
A70.1=Benoni: Klassisk
A70.2=Benoni: Klassisk, 7...a6
A70.3=Benoni: Klassisk, 7...a6 8.a4
A70.4=Benoni: Klassisk, 7...a6 8.a4 Bg4
A70.5=Benoni: Klassisk, 7...a6 8.a4 Bg4 9.Be2
A70.6=Benoni: Klassisk, 7...Bg7
A70.7=Benoni: Klassisk, 8.Be2
A70.8=Benoni: Klassisk, 8.Be2 a6
A70.9=Benoni: Klassisk, 8.Qa4+
A70.10=Benoni: Klassisk, 8.Qa4+ Bd7 9.Qb3 Qc7
A70.11=Benoni: Klassisk, 8.Bf4
A70.12=Benoni: Klassisk, 8.Bf4 O-O 9.Nd2
A70.13=Benoni: Klassisk, 8.Bd3
A70.14=Benoni: Klassisk, 8.Bd3 O-O 9.O-O
A70.15=Benoni: Klassisk, 8.h3
A70.16=Benoni: Klassisk, 8.h3 O-O 9.Bd3
A70.17=Benoni: Klassisk, 8.h3 O-O 9.Bd3 Bd7
A70.18=Benoni: Klassisk, 8.h3 O-O 9.Bd3 Na6
A70.19=Benoni: Klassisk, 8.h3 O-O 9.Bd3 Re8
A70.20=Benoni: Klassisk, 8.h3 O-O 9.Bd3 Re8 10.O-O c4
A70.21=Benoni: Klassisk, 8.h3 O-O 9.Bd3 a6
A70.22=Benoni: Klassisk, 8.h3 O-O 9.Bd3 a6 10.O-O b5
A70.23=Benoni: Klassisk, 8.h3 O-O 9.Bd3 a6 10.a4
A70.24=Benoni: Klassisk, 8.h3 O-O 9.Bd3 a6 10.a4 Nbd7
A70.25=Benoni: Klassisk, 8.h3 O-O 9.Bd3 a6 10.a4 Nbd7 11.O-O Re8
A70.26=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5
A70.27=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5 10.Bxb5
A70.28=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5 10.Nxb5
A70.29=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5 10.Nxb5 Nxe4
A70.30=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5 10.Nxb5 Re8
A70.31=Benoni: Klassisk, 8.h3 O-O 9.Bd3 b5 10.Nxb5 Re8 11.O-O Nxe4
A71.1=Benoni: Klassisk, 8.Bg5
A71.2=Benoni: Klassisk, 8.Bg5 h6 9.Bh4 g5
A71.3=Benoni: Klassisk, 8.Bg5 h6 9.Bh4 a6
A71.4=Benoni: Klassisk, 8.Bg5 h6 9.Bh4 a6 10.Nd2
A71.5=Benoni: Klassisk, 8.Bg5 h6 9.Bh4 a6 10.Nd2 b5 11.Be2
A72.1=Benoni: Klassisk, 8.Be2 O-O
A72.2=Benoni: Klassisk, 8.Be2 O-O 9.Nd2
A72.3=Benoni: Klassisk, 8.Be2 O-O 9.Bg5
A72.4=Benoni: Klassisk, 8.Be2 O-O 9.Bg5 h6 10.Bh4 g5 11.Bg3 Nh5 12.Nd2
A72.5=Benoni: Klassisk, 8.Be2 O-O 9.Bf4
A72.6=Benoni: Klassisk, 8.Be2 O-O 9.Bf4 b5
A72.7=Benoni: Klassisk, 8.Be2 O-O 9.Bf4 a6
A73.1=Benoni: Klassisk, 9.O-O
A73.2=Benoni: Klassisk, 9.O-O Nbd7
A73.3=Benoni: Klassisk, 9.O-O Na6
A73.4=Benoni: Klassisk, 9.O-O Na6 10.Nd2
A73.5=Benoni: Klassisk, 9.O-O Na6 10.Nd2 Nc7
A73.6=Benoni: Klassisk, 9.O-O Bg4
A73.7=Benoni: Klassisk, 9.O-O Bg4 10.Bg5
A73.8=Benoni: Klassisk, 9.O-O Bg4 10.Bf4
A73.9=Benoni: Klassisk, 9.O-O Bg4 10.h3
A73.10=Benoni: Klassisk, 9.O-O a6
A74.1=Benoni: Klassisk, 9.O-O a6 10.a4
A74.2=Benoni: Klassisk, 9.O-O a6 10.a4 Nbd7
A74.3=Benoni: Klassisk, 9.O-O a6 10.a4 Nbd7 11.Nd2
A74.4=Benoni: Klassisk, 9.O-O a6 10.a4 Nbd7 11.Bg5
A74.5=Benoni: Klassisk, 9.O-O a6 10.a4 Nbd7 11.Bf4
A74.6=Benoni: Klassisk, 9.O-O a6 10.a4 Nbd7 11.Bf4 Qe7
A75.1=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4
A75.2=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.h3
A75.3=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Nd2
A75.4=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bg5
A75.5=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bg5 h6
A75.6=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4
A75.7=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Qe7
A75.8=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Re8
A75.9=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Re8 12.Nd2 Bxe2 13.Qxe2 Nh5
A75.10=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Bxf3
A75.11=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Bxf3 12.Bxf3 Qe7
A75.12=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Bxf3 12.Bxf3 Qe7 13.Re1
A75.13=Benoni: Klassisk, 9.O-O a6 10.a4 Bg4 11.Bf4 Bxf3 12.Bxf3 Qe7 med 14.a5
A76.1=Benoni: Klassisk, Huvudvarianten
A76.2=Benoni: Klassisk, Huvudvarianten, 10.Qc2
A76.3=Benoni: Klassisk, Huvudvarianten, 10.Qc2 Bg4
A76.4=Benoni: Klassisk, Huvudvarianten, 10.Qc2 Na6
A76.5=Benoni: Klassisk, Huvudvarianten, 10.Qc2 Na6 11.Bf4
A76.6=Benoni: Klassisk, Huvudvarianten, 10.Qc2 Na6 11.Re1
A76.7=Benoni: Klassisk, Huvudvarianten, 10.Qc2 Na6 11.Re1 Bg4
A77.1=Benoni: Klassisk, Huvudvarianten, 10.Nd2
A77.2=Benoni: Klassisk, Huvudvarianten, 10.Nd2 a6
A77.3=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7
A77.4=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4
A77.5=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 a6
A77.6=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 a6 12.Ra3
A77.7=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 a6 12.Qc2
A77.8=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 a6 12.h3
A77.9=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 Ne5
A77.10=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 Ne5 12.Ndb1
A77.11=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 Ne5 12.Ra3
A77.12=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 Ne5 12.Re1
A77.13=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Nbd7 11.a4 Ne5 12.Qc2
A78.1=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6
A78.2=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.Kh1
A78.3=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.Rb1
A78.4=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.Re1
A79.1=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3
A79.2=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7
A79.3=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7 12.a4
A79.4=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7 12.a4 Nd7
A79.5=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7 12.a4 b6
A79.6=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7 12.a4 b6 13.Kh1
A79.7=Benoni: Klassisk, Huvudvarianten, 10.Nd2 Na6 11.f3 Nc7 12.a4 b6 13.Nc4
A80.1=Holl�ndsk
A80.2=Holl�ndsk: Krejciks gambit
A80.3=Holl�ndsk: Antagen Krejciks gambit
A80.4=Holl�ndsk: Korchnoi attack
A80.5=Holl�ndsk: Korchnoi, Janzen gambit
A80.6=Holl�ndsk: 2.Bg5
A80.7=Holl�ndsk: 2.Bg5 d5
A80.8=Holl�ndsk: 2.Bg5 c6
A80.9=Holl�ndsk: 2.Bg5 Nf6
A80.10=Holl�ndsk: 2.Bg5 h6
A80.11=Holl�ndsk: 2.Bg5 g6
A80.12=Holl�ndsk: 2.Bg5 g6 3.Nc3
A80.13=Holl�ndsk: Alapin
A80.14=Holl�ndsk: Alapin, Manhattan gambit
A80.15=Holl�ndsk: Von Pretzels gambit
A80.16=Holl�ndsk: 2.Nc3
A80.17=Holl�ndsk: 2.Nc3 d5
A80.18=Holl�ndsk: Euwes gambit,2.Nc3 d5 3.e4
A80.19=Holl�ndsk: 2.Nc3 d5 3.Bg5
A80.20=Holl�ndsk: 2.Nc3 Nf6
A80.21=Holl�ndsk: Spielmanns gambit
A80.22=Holl�ndsk: 2.Nc3 Nf6 3.Bg5
A80.23=Holl�ndsk: 2.Nc3 Nf6 3.Bg5 e6
A80.24=Holl�ndsk: 2.Nc3 Nf6 3.Bg5 d5
A80.25=Holl�ndsk: 2.Nc3 Nf6 3.Bg5 d5 4.Bxf6 exf6
A80.26=Holl�ndsk: 2.Nc3 Nf6 3.Bg5 d5 4.Bxf6 exf6 5.e3
A80.27=Holl�ndsk: 2.Nc3 Nf6 3.Bg5 d5 4.Bxf6 exf6 5.e3 c6
A80.28=Holl�ndsk: 2.Nf3
A80.29=Holl�ndsk: 2.Nf3 e6
A80.30=Holl�ndsk: 2.Nf3 e6 3.d5
A80.31=Holl�ndsk: 2.Nf3 Nf6
A80.32=Holl�ndsk: Barczasystemet
A80.33=Holl�ndsk: 2.Nf3 Nf6 3.Bg5
A81.1=Holl�ndsk: 2.g3
A81.2=Holl�ndsk: 2.g3 e6
A81.3=Holl�ndsk: 2.g3 e6 3.Nf3
A81.4=Holl�ndsk: 2.g3 e6 3.Nf3 Nf6
A81.5=Holl�ndsk: 2.g3 Nf6
A81.6=Holl�ndsk: 2.g3 Nf6 3.Nf3
A81.7=Holl�ndsk: 2.g3 Nf6 3.Bg2
A81.8=Holl�ndsk: 2.g3 Nf6 3.Bg2 e6
A81.9=Holl�ndsk: Blackburnevarianten
A81.10=Holl�ndsk: 2.g3 Nf6 3.Bg2 g6
A81.11=Holl�ndsk: 2.g3 Nf6 3.Bg2 g6 4.Nf3
A81.12=Holl�ndsk: Leningrad, Basmanvarianten
A81.13=Holl�ndsk: Leningrad, Carlsbadvarianten
A82.1=Holl�ndsk: Stauntons gambit
A82.2=Holl�ndsk: Stauntons gambit, Baloghs f�rsvar
A82.3=Holl�ndsk: Antagen Stauntons gambit
A82.4=Holl�ndsk: Stauntons gambit, 3.Nc3
A82.5=Holl�ndsk: Stauntons gambit, 3.Nc3 e6
A82.6=Holl�ndsk: Stauntons gambit, 3.Nc3 g6
A82.7=Holl�ndsk: Stauntons gambit, 3.Nc3 Nf6
A82.8=Holl�ndsk: Stauntons gambit, Tartakowervarianten
A82.9=Holl�ndsk: Stauntons gambit, 4.f3
A82.10=Holl�ndsk: Stauntons gambit, 4.f3 e6
A82.11=Holl�ndsk: Stauntons gambit, 4.f3 Nc6
A82.12=Holl�ndsk: Stauntons gambit, 4.f3 exf3
A82.13=Holl�ndsk: Stauntons gambit, 4.f3 exf3 5.Nxf3
A82.14=Holl�ndsk: Stauntons gambit, 4.f3 d5
A82.15=Holl�ndsk: Stauntons gambit, 4.f3 d5 5.fxe4
A83.1=Holl�ndsk: Stauntons gambit, Stauntonvarianten
A83.2=Holl�ndsk: Stauntons gambit, Nimzowitschvarianten
A83.3=Holl�ndsk: Stauntons gambit, Chigorinvarianten
A83.4=Holl�ndsk: Stauntons gambit, 4.Bg5 g6
A83.5=Holl�ndsk: Stauntons gambit, Alekhinevarianten
A83.6=Holl�ndsk: Stauntons gambit, Laskervarianten
A83.7=Holl�ndsk: Stauntons gambit, 4.Bg5 e6
A83.8=Holl�ndsk: Stauntons gambit, 4.Bg5 e6 5.Nxe4
A83.9=Holl�ndsk: Stauntons gambit, 4.Bg5 e6 5.Nxe4 Be7 6.Bxf6 Bxf6 7.Nf3
A83.10=Holl�ndsk: Stauntons gambit, 4.Bg5 Nc6
A83.11=Holl�ndsk: Stauntons gambit, 4.Bg5 Nc6 5.f3
A83.12=Holl�ndsk: Stauntons gambit, 4.Bg5 Nc6 5.d5
A83.13=Holl�ndsk: Stauntons gambit, 4.Bg5 Nc6 5.d5 Ne5 6.Qd4
A84.1=Holl�ndsk: 2.c4
A84.2=Holl�ndsk: 2.c4 d6
A84.3=Holl�ndsk: 2.c4 g6
A84.4=Holl�ndsk: Bladelvarianten
A84.5=Holl�ndsk: 2.c4 e6
A84.6=Holl�ndsk: 2.c4 e6 3.Nf3
A84.7=Holl�ndsk: 2.c4 e6 3.Nf3 Nf6
A84.8=Holl�ndsk: Rubinsteinvarianten
A84.9=Holl�ndsk: Rubinstein, 3...d5
A84.10=Holl�ndsk: Rubinstein, 3...d5 4.e3 c6
A84.11=Holl�ndsk: Avb�jd Stauntons gambit
A84.12=Holl�ndsk: 2.c4 Nf6
A84.13=Holl�ndsk: 2.c4 Nf6 3.Nf3
A85.1=Holl�ndsk: 2.c4 Nf6 3.Nc3
A85.2=Holl�ndsk: 2.c4 Nf6 3.Nc3 d6
A85.3=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6
A85.4=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.a3
A85.5=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.Qc2
A85.6=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.Bg5
A85.7=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.e3
A85.8=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.e3 d5
A85.9=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.e3 Bb4
A85.10=Holl�ndsk: 2.c4 Nf6 3.Nc3 e6 4.Nf3
A85.11=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6
A85.12=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.f3
A85.13=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Bg5
A85.14=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Nf3
A85.15=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Nf3 Bg7
A85.16=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Nf3 Bg7 5.e3
A85.17=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Nf3 Bg7 5.Bf4
A85.18=Holl�ndsk: 2.c4 Nf6 3.Nc3 g6 4.Nf3 Bg7 5.Bg5
A86.1=Holl�ndsk: 2.c4 Nf6 3.g3
A86.2=Holl�ndsk: 2.c4 Nf6 3.g3 d6
A86.3=Holl�ndsk: Hort-Antoshinsystemet
A86.4=Holl�ndsk: Leningradvarianten
A86.5=Holl�ndsk: Leningrad, 4.Nc3
A86.6=Holl�ndsk: Leningrad, 4.Nc3 Bg7
A86.7=Holl�ndsk: Leningrad, 4.Nf3
A86.8=Holl�ndsk: Leningrad, 4.Nf3 Bg7
A86.9=Holl�ndsk: Leningrad, 4.Nf3 Bg7 5.Nc3
A86.10=Holl�ndsk: Leningrad, 4.Bg2
A86.11=Holl�ndsk: Leningrad, 4.Bg2 d6
A86.12=Holl�ndsk: Leningrad, 4.Bg2 Bg7
A86.13=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nh3
A86.14=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3
A86.15=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3 d6
A86.16=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3 d6 6.Nh3
A86.17=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3 d6 6.d5
A86.18=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3 O-O
A86.19=Holl�ndsk: Leningrad, 4.Bg2 Bg7 5.Nc3 O-O 6.Nh3
A87.1=Holl�ndsk: Leningrad, Huvudvarianten
A87.2=Holl�ndsk: Leningrad, Huvudvarianten, 5...d6
A87.3=Holl�ndsk: Leningrad, Huvudvarianten, 5...d6 6.Nc3
A87.4=Holl�ndsk: Leningrad, Huvudvarianten, 5...O-O
A87.5=Holl�ndsk: Leningrad, Huvudvarianten, 6.Nc3
A87.6=Holl�ndsk: Leningrad, Huvudvarianten, 6.Nc3 d6
A87.7=Holl�ndsk: Leningrad, Huvudvarianten, 6.O-O
A87.8=Holl�ndsk: Leningrad, Huvudvarianten, 6...c6
A87.9=Holl�ndsk: Leningrad, Huvudvarianten, 6...d6
A87.10=Holl�ndsk: Leningrad, Huvudvarianten, 7.b3
A87.11=Holl�ndsk: Leningrad, Huvudvarianten, 7.b3 c6
A87.12=Holl�ndsk: Leningrad, Huvudvarianten, 7.d5
A87.13=Holl�ndsk: Leningrad, Huvudvarianten, 7.d5 c6
A87.14=Holl�ndsk: Leningrad, Huvudvarianten, 7.d5 c5
A87.15=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3
A87.16=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 e6
A87.17=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Na6
A87.18=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8
A87.19=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.Re1
A87.20=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.Nd5
A87.21=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.b3
A87.22=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.d5
A87.23=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.d5 a5
A87.24=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.d5 Na6
A87.25=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Qe8 8.d5 Na6 9.Rb1
A88.1=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6
A88.2=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.Re1
A88.3=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.Qc2
A88.4=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.b3
A88.5=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.b3 Na6
A88.6=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.b3 Qe8
A88.7=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.b3 Qa5
A88.8=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5
A88.9=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 cxd5
A88.10=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 Qe8
A88.11=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 Qa5
A88.12=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 Bd7
A88.13=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 e5
A88.14=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 e5 9.dxe6 Bxe6 10.b3
A88.15=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 c6 8.d5 e5 9.dxe6 Bxe6 10.Qd3
A89.1=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6
A89.2=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.b3
A89.3=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5
A89.4=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Na5
A89.5=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Na5 9.Qd3
A89.6=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Na5 9.Nd2
A89.7=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Ne5
A89.8=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Ne5 9.Nxe5
A89.9=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Ne5 9.Nxe5 dxe5 10.Qb3
A89.10=Holl�ndsk: Leningrad, Huvudvarianten, 7.Nc3 Nc6 8.d5 Ne5 9.Nxe5 dxe5 10.e4
A90.6=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2
A90.7=Holl�ndsk: Holl�ndsk-Indisk (Nimzo-Holl�ndsk)varianten
A90.8=Holl�ndsk: Holl�ndsk-Indisk, 5.Nc3
A90.9=Holl�ndsk: Holl�ndsk-Indisk, 5.Nd2
A90.10=Holl�ndsk: Holl�ndsk-Indisk, 5.Bd2
A90.11=Holl�ndsk: Holl�ndsk-Indisk, Alekhinevarianten
A90.12=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 d5
A90.13=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 d5 5.Nh3
A90.14=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 d5 5.Nf3
A90.15=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 c6
A90.16=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 c6 5.Nh3
A90.17=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 c6 5.Nf3
A90.18=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 c6 5.Nf3 d5
A90.19=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.Nc3
A90.20=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.Qc2
A90.21=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.Qc2 Bd6
A90.22=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.O-O
A90.23=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.O-O Bd6
A90.24=Holl�ndsk: 2.c4 Nf6 3.g3 e6 5.Nf3 d5 6.O-O Bd6 7.b3
A91.1=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7
A91.2=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3
A91.3=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3 O-O 6.O-O
A91.4=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3 O-O 6.O-O d6
A91.5=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3 O-O 6.O-O d6 7.Nc3
A91.6=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3 O-O 6.O-O d6 7.Nc3 c6
A91.7=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nh3 O-O 6.O-O d6 7.Nc3 Qe8
A91.8=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nc3
A91.9=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nc3 d5
A91.10=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nc3 O-O
A91.11=Holl�ndsk: Botvinnik-Bronsteinvarianten, 5.Nc3 O-O 6.e3
A91.12=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3
A91.13=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 d6
A91.14=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 d6 6.Nc3
A91.15=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 d5
A91.16=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 d5 6.O-O
A91.17=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 d5 6.O-O c6
A92.1=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O
A92.2=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.d5
A92.3=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.Nc3
A92.4=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.Nc3 d6
A92.5=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.O-O
A92.6=Holl�ndsk: Alekhinevarianten
A92.7=Holl�ndsk: Alekhine, 7.d5
A92.8=Holl�ndsk: Alekhine, 7.Nbd2
A92.9=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.O-O c6
A92.10=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.O-O c6 7.b3
A92.11=Holl�ndsk: 2.c4 Nf6 3.g3 e6 4.Bg2 Be7 5.Nf3 O-O 6.O-O c6 7.b3 a5
A92.12=Holl�ndsk: Stonewallvarianten
A92.13=Holl�ndsk: Stonewall, 7.Nbd2
A92.14=Holl�ndsk: Stonewall, 7.Nbd2 c6
A92.15=Holl�ndsk: Stonewall, 7.Qc2
A92.16=Holl�ndsk: Stonewall, 7.Qc2 c6
A92.17=Holl�ndsk: Stonewall, 7.Qc2 c6 8.Nbd2
A92.18=Holl�ndsk: Stonewall, 7.Nc3
A93.1=Holl�ndsk: Stonewall, Botvinnikvarianten
A93.2=Holl�ndsk: Stonewall, Botvinnik, 7...b6
A93.3=Holl�ndsk: Stonewall, Botvinnik, 7...Nc6
A93.4=Holl�ndsk: Stonewall, Botvinnik, 7...c6
A93.5=Holl�ndsk: Stonewall, Botvinnik, 8.Bb2
A93.6=Holl�ndsk: Stonewall, Botvinnik, 8.Qc2
A93.7=Holl�ndsk: Stonewall, Botvinnik, 8.Qc2 Ne4
A94.1=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3
A94.2=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bd7
A94.3=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Nbd7
A94.4=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Nbd7 9.Bxe7
A94.5=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bxa3
A94.6=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bxa3 9.Nxa3
A94.7=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bxa3 9.Nxa3 Nbd7
A94.8=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bxa3 9.Nxa3 Qe7
A94.9=Holl�ndsk: Stonewall, Botvinnik, 8.Ba3 Bxa3 9.Nxa3 Qe7 10.Qc1
A95.1=Holl�ndsk: Stonewall, 7.Nc3 c6
A95.2=Holl�ndsk: Stonewall, 7.Nc3 c6 8.Ne5
A95.3=Holl�ndsk: Stonewall, 7.Nc3 c6 8.Bf4
A95.4=Holl�ndsk: Stonewall, 7.Nc3 c6 8.Bg5
A95.5=Holl�ndsk: Stonewall, 7.Nc3 c6 8.Qc2
A95.6=Holl�ndsk: Stonewall: Chekhovervarianten, 8.Qc2 Qe8 9.Bg5
A95.7=Holl�ndsk: Stonewall, 7.Nc3 c6 8.b3
A95.8=Holl�ndsk: Stonewall, 7.Nc3 c6 8.b3 Qe8
A96.1=Holl�ndsk: Klassisk
A96.2=Holl�ndsk: Klassisk, 7.b3
A96.3=Holl�ndsk: Klassisk, 7.b3 a5
A96.4=Holl�ndsk: Klassisk, 7.b3 a5 8.Bb2
A96.5=Holl�ndsk: Klassisk, 7.b3 Qe8
A96.6=Holl�ndsk: Klassisk, 7.b3 Qe8 8.Bb2
A96.7=Holl�ndsk: Klassisk, 7.Nc3
A96.8=Holl�ndsk: Klassisk, 7.Nc3 a5
A96.9=Holl�ndsk: Klassisk, 7.Nc3 a5 8.Qc2
A96.10=Holl�ndsk: Klassisk, 7.Nc3 a5 8.Re1
A96.11=Holl�ndsk: Klassisk, 7.Nc3 a5 8.b3
A97.1=Holl�ndsk: Ilyin-Zhenevskyvarianten
A97.2=Holl�ndsk: Ilyin-Zhenevsky, 8.b4
A97.3=Holl�ndsk: Ilyin-Zhenevsky, Wintervarianten
A97.4=Holl�ndsk: Ilyin-Zhenevsky, Winter, 8...Ne4
A97.5=Holl�ndsk: Ilyin-Zhenevsky, Winter, 8...Qg6
A97.6=Holl�ndsk: Ilyin-Zhenevsky, Winter, 8...Qg6 9.e4
A98.1=Holl�ndsk: Ilyin-Zhenevsky, 8.Qc2
A98.2=Holl�ndsk: Ilyin-Zhenevsky, 8.Qc2 Nc6
A98.3=Holl�ndsk: Ilyin-Zhenevsky, 8.Qc2 Qh5
A99.1=Holl�ndsk: Ilyin-Zhenevsky, 8.b3
A99.2=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 Qh5
A99.3=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 a5
A99.4=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 a5 9.Qc2
A99.5=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 a5 9.Bb2
A99.6=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 a5 9.Bb2 Na6
A99.7=Holl�ndsk: Ilyin-Zhenevsky, 8.b3 a5 9.Bb2 Qh5
B00.1=Kungsbondespel
B00.2=Kungsbonde: Flodh�stf�rsvaret
B00.3=Kungsbonde: Fred
B00.4=Omv�nd Grob (Borg/Basman-f�rsvaret)
B00.5=Omv�nd Grob (Borg/Basman-f�rsvaret)
B00.6=St. Georges f�rsvar
B00.7=St. Georges f�rsvar
B00.8=Hemsk krypande omv�nd (Basman) �ppning
B00.9=Owens f�rsvar
B00.10=Owens f�rsvar
B00.11=Owens f�rsvar: Fransk
B00.12=Owens f�rsvar: 2.d4 Bb7
B00.13=Owens f�rsvar: Naselwaus gambit
B00.14=Owens f�rsvar: Smiths gambit
B00.15=Owens f�rsvar: 3.Bd3
B00.16=Owens f�rsvar: Matinovskys gambit
B00.17=Owens f�rsvar: 3.Bd3 Nf6
B00.18=Owens f�rsvar: 3.Bd3 e6
B00.19=Owens f�rsvar: 3.Bd3 e6 4.Nf3
B00.20=Owens f�rsvar: 3.Bd3 e6 4.Nf3 c5
B00.21=Owens f�rsvar: 3.Bd3 e6 4.Nf3 c5 5.c3
B00.22=Nimzowitsch f�rsvar
B00.23=Nimzowitsch f�rsvar: Wheelers gambit
B00.24=Nimzowitsch f�rsvar: 2.Nc3
B00.25=Nimzowitsch f�rsvar: 2.Nc3 e6
B00.26=Nimzowitsch f�rsvar: 2.Nf3
B00.27=Nimzowitsch f�rsvar: Colorados motangrepp
B00.28=Nimzowitsch f�rsvar: 2.Nf3 d6
B00.29=Nimzowitsch f�rsvar: 2.Nf3 d6 3.d4 Nf6
B00.30=Nimzowitsch f�rsvar: 2.Nf3 d6 3.d4 Nf6 4.Nc3
B00.31=Nimzowitsch f�rsvar: 2.Nf3 d6 3.d4 Nf6 4.Nc3 Bg4
B00.32=Nimzowitsch f�rsvar: 2.Nf3 d6 3.d4 Nf6 4.Nc3 Bg4 5.Be2
B00.33=Nimzowitsch f�rsvar: 2.Nf3 d6 3.d4 Nf6 4.Nc3 Bg4 5.Be3
B00.34=Nimzowitsch f�rsvar: 2.d4
B00.35=Nimzowitsch f�rsvar: 2.d4 e5
B00.36=Nimzowitsch f�rsvar: 2.d4 e5 3.dxe5
B00.37=Nimzowitsch f�rsvar: Bielefelders gambit
B00.38=Nimzowitsch f�rsvar: 2.d4 e5 3.d5
B00.39=Nimzowitsch f�rsvar: 2.d4 d5
B00.40=Nimzowitsch f�rsvar: 2.d4 d5 3.exd5
B00.41=Nimzowitsch f�rsvar: Aachens gambit
B00.42=Nimzowitsch f�rsvar: 2.d4 d5 3.exd5 Qxd5
B00.43=Nimzowitsch f�rsvar: Marshalls gambit
B00.44=Nimzowitsch f�rsvar: 2.d4 d5 3.exd5 Qxd5 4.Nf3
B00.45=Nimzowitsch f�rsvar: Bogoljubowvarianten
B00.46=Nimzowitsch f�rsvar: Bogoljubow, 3...dxe4
B00.47=Nimzowitsch f�rsvar: 2.d4 d5 3.e5
B01.1=Skandinavisk (Centrummotangepp)
B01.2=Skandinavisk: 2.d3
B01.3=Skandinavisk: 2.e5
B01.4=Skandinavisk: 2.exd5
B01.5=Skandinavisk: B�hnkes gambit
B01.6=Skandinavisk: 2...Qxd5
B01.7=Skandinavisk: 2...Qxd5 3.Nf3
B01.8=Skandinavisk: 2...Qxd5 3.Nf3 Nf6
B01.9=Skandinavisk: 2...Qxd5 3.d4
B01.10=Skandinavisk: 2...Qxd5 3.d4 Nf6
B01.11=Skandinavisk: 2...Qxd5 3.d4 e5
B01.12=Skandinavisk: 2...Qxd5 3.Nc3
B01.13=Skandinavisk: 2...Qxd5 3.Nc3 Qd8
B01.14=Skandinavisk: Schillers f�rsvar
B01.15=Skandinavisk: Schiller, 4.d4 Nf6
B01.16=Skandinavisk: Schiller, Bronsteinvarianten
B01.17=Skandinavisk: 2...Qxd5 3.Nc3 Qa5
B01.18=Skandinavisk, Mieses gambit
B01.19=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.g3
B01.20=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.Bc4
B01.21=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.Bc4 Nf6
B01.22=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.Nf3
B01.23=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.Nf3 Nf6
B01.24=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.Nf3 Nf6 5.Be2
B01.25=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.d4
B01.26=Skandinavisk: Anderssens motattack
B01.27=Skandinavisk: Anderssens motattack, G�teborgsvarianten
B01.28=Skandinavisk: Anderssens motattack, Collijnvarianten
B01.29=Skandinavisk: Anderssens motattack, 5.dxe5
B01.30=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.d4 c6
B01.31=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.d4 c6 5.Bc4
B01.32=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.d4 c6 5.Nf3
B01.33=Skandinavisk: 2...Qxd5 3.Nc3 Qa5 4.d4 Nf6
B01.34=Skandinavisk: 2...Qxd5, 5.Bd2
B01.35=Skandinavisk: 2...Qxd5, 5.Bd2 c6
B01.36=Skandinavisk: 2...Qxd5, 5.Bc4
B01.37=Skandinavisk: 2...Qxd5, 5.Bc4 c6
B01.38=Skandinavisk: 2...Qxd5, 5.Nf3
B01.39=Skandinavisk: 2...Qxd5, 5.Nf3 Bg4
B01.40=Skandinavisk: Laskervarianten
B01.41=Skandinavisk: 2...Qxd5, 5.Nf3 Bf5
B01.42=Skandinavisk: Gr�nfeldvarianten
B01.43=Skandinavisk: 2...Qxd5, 5.Nf3 Bf5 6.Bc4
B01.44=Skandinavisk: 2...Qxd5, Huvudvarianten
B01.45=Skandinavisk: 2...Qxd5, Huvudvarianten, 6.Bc4
B01.46=Skandinavisk: 2...Qxd5, Huvudvarianten, 6.Bc4 Bg4
B01.47=Skandinavisk: 2...Qxd5, Huvudvarianten, 6.Bc4 Bf5
B01.48=Skandinavisk: 2...Qxd5, Huvudvarianten, 6.Bc4 Bf5 7.Bd2
B01.49=Skandinavisk: 2...Qxd5, Huvudvarianten, 6.Bc4 Bf5 7.Bd2 e6
B01.50=Skandinavisk: 2...Qxd5, Huvudvarianten, 8.Nd5
B01.51=Skandinavisk: 2...Qxd5, Huvudvarianten, 8.Qe2
B01.52=Skandinavisk: 2...Qxd5, Huvudvarianten, 8.Qe2 Bb4
B01.53=Skandinavisk: 2...Qxd5, Huvudvarianten, 8.Qe2 Bb4 9.a3
B01.54=Skandinavisk: 2...Qxd5, Huvudvarianten, 8.Qe2 Bb4 9.O-O-O
B01.55=Skandinavisk: 2...Nf6
B01.56=Skandinavisk: 2...Nf6 3.Bc4
B01.57=Skandinavisk: 2...Nf6 3.Nf3
B01.58=Skandinavisk: 2...Nf6 3.Nf3 Nxd5
B01.59=Skandinavisk: 2...Nf6 3.Bb5+
B01.60=Skandinavisk: 2...Nf6 3.Bb5+ Nbd7
B01.61=Skandinavisk: 2...Nf6 3.Bb5+ Bd7
B01.62=Skandinavisk: 2...Nf6 3.Bb5+ Bd7 4.Bc4
B01.63=Skandinavisk: 2...Nf6 3.Bb5+ Bd7 4.Bc4 Bg4
B01.64=Skandinavisk: 2...Nf6 3.Bb5+ Bd7 4.Be2
B01.65=Skandinavisk: 2...Nf6 3.Bb5+ Bd7 4.Be2 Nxd5 5.d4 Bf5
B01.66=Skandinavisk: 2...Nf6 3.c4
B01.67=Skandinavisk: Skandinavisk gambit
B01.68=Skandinavisk: Antagen Skandinavisk gambit
B01.69=Skandinavisk: Isl�ndsk gambit
B01.70=Skandinavisk: Antagen Isl�ndsk gambit, 4.dxe6
B01.71=Skandinavisk: Antagen Isl�ndsk gambit, 4.dxe6 Bxe6
B01.72=Skandinavisk: Antagen Isl�ndsk gambit, 4.dxe6 Bxe6 5.d4
B01.73=Skandinavisk: Antagen Isl�ndsk gambit, 4.dxe6 Bxe6 5.Nf3
B01.74=Skandinavisk: 2...Nf6 3.d4
B01.75=Skandinavisk: Richtervarianten
B01.76=Skandinavisk: Portuguisiska varianten
B01.77=Skandinavisk: Portuguisiska, 4.Bb5+
B01.78=Skandinavisk: Portuguisiska, 4.Nf3
B01.79=Skandinavisk: Portuguisiska, 4.Nf3 Qxd5
B01.80=Skandinavisk: Portuguisiska, 4.Nf3 Qxd5 5.Be2
B01.81=Skandinavisk: Portuguisiska, 4.Nf3 Qxd5 5.Be2 Nc6
B01.82=Skandinavisk: Portuguisiska, 4.Be2
B01.83=Skandinavisk: Portuguisiska, 4.Be2 Bxe2
B01.84=Skandinavisk: Portuguisiska, 4.f3
B01.85=Skandinavisk: Portuguisiska, 4.f3 Bf5
B01.86=Skandinavisk: Portuguisiska, 4.f3 Bf5 5.c4
B01.87=Skandinavisk: Portuguisiska, 4.f3 Bf5 5.Bb5+
B01.88=Skandinavisk: Portuguisiska, 4.f3 Bf5 5.Bb5+ Nbd7
B01.89=Skandinavisk: Portuguisiska, 4.f3 Bf5 5.Bb5+ Nbd7 6.c4
B01.90=Skandinavisk: Marshallvarianten
B01.91=Skandinavisk: Marshall, 4.Nf3
B01.92=Skandinavisk: Marshall, 4.Nf3 Bf5
B01.93=Skandinavisk: Marshall, 4.Nf3 Bg4
B01.94=Skandinavisk: Marshall, 4.Nf3 Bg4 5.Be2
B01.95=Skandinavisk: Marshall, 4.Nf3 Bg4 5.Be2 e6
B01.96=Skandinavisk: Marshall, 4.Nf3 g6
B01.97=Skandinavisk: Marshall, 4.Nf3 g6 5.Be2
B01.98=Skandinavisk: Marshall, 4.Nf3 g6 5.Be2 Bg7
B01.99=Skandinavisk: Marshall, 4.c4
B01.10=Skandinavisk: Marshall, 4.c4 Nf6
B01.10=Skandinavisk: Marshall, 4.c4 Nb6
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nc3
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nc3 e5
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 Bg4
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 Bg4 6.Be2 e6
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 Bg4 6.c5
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6
B01.10=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.Be2
B01.11=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.Be2 Bg7
B01.11=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.h3
B01.11=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.h3 Bg7
B01.11=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.Nc3
B01.11=Skandinavisk: Marshall, 4.c4 Nb6 5.Nf3 g6 6.Nc3 Bg7
B02.1=Alekhines f�rsvar
B02.2=Alekhine: Krejcikvarianten
B02.3=Alekhine: Maroczyvarianten
B02.4=Alekhine: Skandinavisk variant
B02.5=Alekhine: Skandinavisk variant, 2.Nc3 d5
B02.6=Alekhine: Skandinavisk, 3.e5
B02.7=Alekhine: Skandinavisk, 3.e5 Ne4
B02.8=Alekhine: Skandinavisk, 3.e5 Nfd7
B02.9=Alekhine: Spielmanns gambit
B02.10=Alekhine: Skandinavisk, Avbyte
B02.11=Alekhine: Skandinavisk, Geschevs gambit
B02.12=Alekhine: Skandinavisk, Avbyte
B02.13=Alekhine: Skandinavisk, Avbyte, 4.Nf3
B02.14=Alekhine: Skandinavisk, Avbyte, 4.Nxd5
B02.15=Alekhine: Skandinavisk, Avbyte, 4.Nxd5
B02.16=Alekhine: Skandinavisk, Avbyte, 4.Bc4
B02.17=Alekhine: Skandinavisk, Avbyte, 4.Bc4 Nb6
B02.18=Alekhine: 2.e5
B02.19=Alekhine: Mokele Mbembe (B�cker)varianten
B02.20=Alekhine: Brooklyns f�rsvar (Retr�ttvarianten)
B02.21=Alekhine: 2.e5 Nd5
B02.22=Alekhine: Wellingvarianten
B02.23=Alekhine: 3.Bc4
B02.24=Alekhine: Kmochvarianten
B02.25=Alekhine: S�misch attack
B02.26=Alekhine: S�misch attack, 3...Nxc3
B02.27=Alekhine: Chasevarianten
B02.28=Alekhine: Chasevarianten, 3.c4 Nb6
B02.29=Alekhine: Chase, Steinervarianten
B02.30=Alekhine: Tv�bonde (Lasker) attack
B02.31=Alekhine: Tv�bondeattack, 5.Nc3
B02.32=Alekhine: Tv�bondeattack, 5.Bc4
B02.33=Alekhine: Tv�bondeattack, Mikenasvarianten
B03.1=Alekhine: 3.d4
B03.2=Alekhine: O'Sullivans gambit
B03.3=Alekhine: 3.d4 d6
B03.4=Alekhine: 3.d4 d6 4.exd6
B03.5=Alekhine: Baloghvarianten, 1.e4 Nf6 2.e5 Nd5 3.d4 d6 4.Bc4
B03.6=Alekhine: 4.c4
B03.7=Alekhine: 4.c4 Nb6
B03.8=Alekhine: 4.c4 Nb6 5.Nf3
B03.9=Alekhine: Fyrbondeattack
B03.10=Alekhine: Fyrbondeattack, Planincvarianten
B03.11=Alekhine: Fyrbondeattack, Trifunovicvarianten
B03.12=Alekhine: Fyrbondeattack, Fianchettovarianten
B03.13=Alekhine: Fyrbondeattack, 5...dxe5
B03.14=Alekhine: Fyrbondeattack, 5...dxe5 6.fxe5
B03.15=Alekhine: Fyrbondeattack, 6...c5
B03.16=Alekhine: Fyrbondeattack, 6...Bf5
B03.17=Alekhine: Fyrbondeattack, Fahrnivarianten
B03.18=Alekhine: Fyrbondeattack, Korchnoivarianten
B03.19=Alekhine: Fyrbondeattack, 6...Nc6
B03.20=Alekhine: Fyrbondeattack, Ilyin-Zhenevskyvarianten
B03.21=Alekhine: Fyrbondeattack, 7.Be3
B03.22=Alekhine: Avbytesvarianten
B03.23=Alekhine: Avbyte, 5...exd6
B03.24=Alekhine: Avbyte, 5...exd6 6.Nc3
B03.25=Alekhine: Avbyte, 5...exd6 6.Nc3 Be7
B03.26=Alekhine: Avbyte, 5...cxd6
B03.27=Alekhine: Avbyte, 5...cxd6 6.Nc3
B03.28=Alekhine: Avbyte, 5...cxd6 6.Nc3 g6 7.Be3
B04.1=Alekhine: Moderna varianten
B04.2=Alekhine: Modern, 4...Nc6
B04.3=Alekhine: Modern, 4...c6
B04.4=Alekhine: Modern, 4...c6 5.c4
B04.5=Alekhine: Modern, Schmidvarianten
B04.6=Alekhine: Modern, Larsenvarianten
B04.7=Alekhine: Modern, Larsen, 5.Nxe5 g6
B04.8=Alekhine: Modern, Larsen, 5.Nxe5 g6 6.Bc4
B04.9=Alekhine: Modern, Larsen, 5.Nxe5 g6 6.Bc4 c6 7.O-O
B04.10=Alekhine: Modern, Fianchettovarianten
B04.11=Alekhine: Modern, Fianchetto, 5.Bc4
B04.12=Alekhine: Modern, Fianchetto, 5.Bc4 Nb6
B04.13=Alekhine: Modern, Fianchetto, 5.Bc4 Nb6 6.Bb3 Bg7
B04.14=Alekhine: Modern, Fianchetto, Keresvarianten
B04.15=Alekhine: Modern, Fianchetto, 5.Bc4 Nb6 6.Bb3 Bg7 7.Ng5
B05.1=Alekhine: Modern, 4...Bg4
B05.2=Alekhine: Modern, Panovvarianten
B05.3=Alekhine: Modern, Alekhinevarianten
B05.4=Alekhine: Modern, Alekhinevarianten, 5.c4 Nb6
B05.5=Alekhine: Modern, Alekhinevarianten, 6.exd6
B05.6=Alekhine: Modern, Alekhinevarianten, 6.exd6 cxd6
B05.7=Alekhine: Modern, Alekhinevarianten, 6.exd6 exd6
B05.8=Alekhine: Modern, 5.Be2
B05.9=Alekhine: Modern, 5.Be2 Nc6
B05.10=Alekhine: Modern, Flohrvarianten
B05.11=Alekhine: Modern, Flohrvarianten, 6.c4
B05.12=Alekhine: Modern, Flohrvarianten, 6.O-O
B05.13=Alekhine: Modern, 5.Be2 e6
B05.14=Alekhine: Modern, 5.Be2 e6 6.O-O
B05.15=Alekhine: Modern, Huvudvarianten
B05.16=Alekhine: Modern, Huvudvarianten, 8.h3
B05.17=Alekhine: Modern, Huvudvarianten, 8.h3 Bh5
B05.18=Alekhine: Modern, Huvudvarianten, 8.h3 Bh5 9.Nc3
B05.19=Alekhine: Modern, Huvudvarianten, 8.h3 Bh5 9.Nc3 O-O
B05.20=Alekhine: Modern, Huvudvarianten, 8.h3 Bh5 9.Nc3 O-O 10.Be3
B05.21=Alekhine: Modern, Huvudvarianten, 8.h3 Bh5 9.Nc3 O-O 10.Be3 d5
B05.22=Alekhine: Modern, Huvudvarianten, 8.exd6
B05.23=Alekhine: Modern, Huvudvarianten, 8.Nc3
B05.24=Alekhine: Modern, Huvudvarianten, 8.Nc3 O-O 9.Be3
B05.25=Alekhine: Modern, Huvudvarianten, 8.Nc3 O-O 9.Be3 Nc6
B05.26=Alekhine: Modern, Huvudvarianten, 8.Nc3 O-O 9.Be3 Nc6 10.exd6 cxd6
B06.1=Modern: 1.e4 g6
B06.2=Modern: 1.e4 g6 2.Nc3
B06.3=Modern: 1.e4 g6 2.Nc3 d6
B06.4=Modern: 1.e4 g6 2.Nc3 Bg7
B06.5=Modern: 1.e4 g6 2.Nc3 Bg7 3.f4 d6
B06.6=Modern: 1.e4 g6 2.f4
B06.7=Modern: 1.e4 g6 2.f4 d6
B06.8=Modern: 1.e4 g6 2.f4 Bg7 3.Nf3
B06.9=Modern: 1.e4 g6 2.f4 Bg7 3.Nf3 d6
B06.10=Modern: 1.e4 g6 2.d4
B06.11=Modern: Norskt f�rsvar
B06.12=Modern: Norskt f�rsvar, 3.e5 Nh5 4.g4 Ng7
B06.13=Modern: 1.e4 g6 2.d4 c6
B06.14=Modern: 1.e4 g6 2.d4 d6
B06.15=Modern: 1.e4 g6 2.d4 Bg7
B06.16=Modern: 1.e4 g6 2.d4 Bg7 3.Bc4
B06.17=Modern: 1.e4 g6 2.d4 Bg7 3.c3
B06.18=Modern: 1.e4 g6 2.d4 Bg7 3.c3 d63.c3
B06.19=Modern: Pterodactyl med c3
B06.20=Modern: Gellersystemet
B06.21=Modern: 3.Nf3
B06.22=Modern: 3.Nf3 d6
B06.23=Modern: 3.Nf3 d6 4.Bc4
B06.24=Modern: 3.Nc3
B06.25=Modern: Mittenbergers gambit
B06.26=Modern: Pterodactyl med Nc3
B06.27=Modern: 3.Nc3
B06.28=Modern: 3.Nc3 d6 4.Bc4
B06.29=Modern: 3.Nc3 d6 4.Bc4 c6
B06.30=Modern: 3.Nc3 d6 4.Bc4 c6 5.Qf3
B06.31=Modern: 3.Nc3 d6 4.Bc4 c6 5.Qf3 Nf6
B06.32=Modern: 3.Nc3 d6 4.Bc4 c6 5.Qf3 e6
B06.33=Modern: 3.Nc3 d6 4.Be3
B06.34=Modern: 3.Nc3 d6 4.Be3 a6
B06.35=Modern: 3.Nc3 d6 4.Be3 c6
B06.36=Modern: Tv� springare-varianten
B06.37=Modern: Tv� springare, Suttlesvarianten
B06.38=Modern: Tv� springare, Suttles, Tal gambit
B06.39=Modern: Pseudo-�sterrikisk attack, 1.e4 g6 2.d4 Bg7 3.Nc3 d6 4.f4
B06.40=Modern: Pseudo-�sterrikisk attack, 1.e4 g6 2.d4 Bg7 3.Nc3 d6 4.f4 c6
B06.41=Modern: Pseudo-�sterrikisk attack, 1.e4 g6 2.d4 Bg7 3.Nc3 d6 4.f4 c6 5.Nf3
B06.42=Modern: Pseudo-�sterrikisk attack, 1.e4 g6 2.d4 Bg7 3.Nc3 d6 4.f4 Nc6
B06.43=Modern: Trebondeattack, 1.e4 g6 2.d4 Bg7 3.f4
B07.1=Pirc: 1.e4 d6
B07.2=Pirc: 1.e4 d6 2.g3
B07.3=Pirc: 1.e4 d6 2.c4
B07.4=Pirc: 2.Nc3
B07.5=Pirc: 2.Nc3 Nf6
B07.6=Pirc: 2.Nf3
B07.7=Pirc-Retis: Wades f�rsvar, 1.e4 d6 2.Nf3 Bg4
B07.8=Pirc: 2.Nf3 Nf6
B07.9=Pirc: 2.Nf3 Nf6 3.Nc3
B07.10=Pirc: 2.f4
B07.11=Pirc: 2.f4 Nf6
B07.12=Pirc: 2.f4 Nf6 3.Nc3
B07.13=Pirc: 2.f4 Nf6 3.Nc3 g6 4.Nf3 Bg7
B07.14=Pirc: 2.d4
B07.15=Pirc: 2.d4 c6
B07.16=Pirc: Lengfellnersystemet
B07.17=Pirc: 2.d4 Nd7
B07.18=Pirc: 2.d4 Nf6
B07.19=Pirc: Roschers gambit
B07.20=Pirc: 3.Nbd2
B07.21=Pirc: 3.Nbd2 g6
B07.22=Pirc: 3.Nbd2 g6
B07.23=Pirc: 3.f3
B07.24=Pirc: 3.f3 e5
B07.25=Pirc: 3.f3 e5 Dambyte
B07.26=Pirc: 3.f3 e5 4.d5
B07.27=Pirc: 3.f3 g6
B07.28=Pirc: 3.Bd3
B07.29=Pirc: 3.Bd3 e5
B07.30=Pirc: 3.Bd3 e5 4.c3 d5
B07.31=Pirc: 3.Bd3 e5 4.c3 d5 5.dxe5 dxe4
B07.32=Pirc: 3.Bd3 e5 4.c3 d5 5.dxe5 Nxe4
B07.33=Pirc: 3.Bd3 g6
B07.34=Pirc: 3.Bd3 g6 4.Nf3
B07.35=Pirc: 3.Bd3 g6 4.Nf3 Bg7
B07.36=Pirc: 3.Bd3 g6 4.Nf3 Bg7 5.c3
B07.37=Pirc: 3.Nc3
B07.38=Pirc: 3.Nc3 Nbd7
B07.39=Pirc: 3.Nc3 e5
B07.40=Pirc: 3.Nc3 e5 Dambyte
B07.41=Pirc: Pytel-Tjeckiskt
B07.42=Pirc: Pytel-Tjeckiskt, 4.Nf3
B07.43=Pirc: Pytel-Tjeckiskt, 4.f4
B07.44=Pirc: Pytel-Tjeckiskt, 4.f4 Qa5
B07.45=Pirc: 3...g6
B07.46=Pirc: 3...g6 4.h4
B07.47=Pirc: 4.Nge2
B07.48=Pirc: 4.Nge2 Bg7
B07.49=Pirc: Sveshnikov, 4.g3
B07.50=Pirc: Sveshnikov, 4.g3 Bg7
B07.51=Pirc: Sveshnikov, 4.g3 Bg7 5.Bg2 c6
B07.52=Pirc: Holmov, 4.Bc4
B07.53=Pirc: Holmov, 4.Bc4 Bg7
B07.54=Pirc: 4.Be3
B07.55=Pirc: 4.Be3 c6
B07.56=Pirc: 4.Be3 Bg7
B07.57=Pirc: 150 attack, 4.Be3 Bg7 5.Qd2
B07.58=Pirc: 150 attack, 4.Be3 Bg7 5.Qd2 c6
B07.59=Pirc: 150 attack, 4.Be3 Bg7 5.Qd2 c6 6.f3 b5
B07.60=Pirc: Byrne 4.Bg5
B07.61=Pirc: 4.Bg5 Bg7
B07.62=Pirc: 4.Be2
B07.63=Pirc: 4.Be2 Bg7
B07.64=Pirc: Kinesiska varianten, 1.e4 d6 2.d4 Nf6 3.Nc3 g6 4.Be2 Bg7 5.g4
B07.65=Pirc: Barjonett-Mariotti attack, 1.e4 d6 2.d4 Nf6 3.Nc3 g6 4.Be2 Bg7 5.h4
B08.1=Pirc: Klassisk, 1.e4 d6 2.d4 Nf6 3.Nc3 g6 4.Nf3
B08.2=Pirc: Klassisk, 4.Nf3 Bg7
B08.3=Pirc: Klassisk, 4.Nf3 Bg7 5.h3
B08.4=Pirc: Klassisk, 4.Nf3 Bg7 5.h3 c6
B08.5=Pirc: Klassisk, 4.Nf3 Bg7 5.h3 O-O
B08.6=Pirc: Klassisk, Spasskysystemet, 1.e4 d6 2.d4 Nf6 3.Nc3 g6 4.Nf3 Bg7 5.h3 O-O 6.Be3
B08.7=Pirc: Klassisk, Spasskysystemet, 6...d5
B08.8=Pirc: Klassisk, Spasskysystemet, 6...a6
B08.9=Pirc: Klassisk, Spasskysystemet, 6...c6
B08.10=Pirc: Klassisk, 5.a4
B08.11=Pirc: Klassisk, 5.a4 c6
B08.12=Pirc: Klassisk, 5.Bc4
B08.13=Pirc: Klassisk, 5.Bc4 c6
B08.14=Pirc: Klassisk, 5.Be3
B08.15=Pirc: Klassisk, 5.Be3 a6 6.a4
B08.16=Pirc: Klassisk, 5.Be3 c6
B08.17=Pirc: Klassisk, 5.Be2
B08.18=Pirc: Klassisk, 5.Be2 a6 6.a4
B08.19=Pirc: Klassisk, 5.Be2 c6
B08.20=Pirc: Klassisk, 5.Be2 O-O
B08.21=Pirc: Klassisk, 5.Be2 O-O 6.Be3
B08.22=Pirc: Klassisk, 5.Be2 O-O 6.O-O
B08.23=Pirc: Klassisk, 5.Be2 O-O 6.O-O Nc6
B08.24=Pirc: Klassisk, 5.Be2 O-O 6.O-O c6
B08.25=Pirc: Klassisk, 5.Be2 O-O 6.O-O c6 7.h3
B08.26=Pirc: Klassisk, 5.Be2 O-O 6.O-O c6 7.a4
B08.27=Pirc: Klassisk, 5.Be2 O-O 6.O-O c6 7.a4 Nbd7
B08.28=Pirc: Klassisk, 5.Be2 O-O 6.O-O Bg4
B08.29=Pirc: Klassisk, 5.Be2 O-O 6.O-O Bg4 7.Be3 Nc6 8.Qd2
B08.30=Pirc: Klassisk, 5.Be2 O-O 6.O-O Bg4 7.Be3 Nc6 8.Qd2 e5
B09.1=Pirc: �sterrikisk attack, 1.e4 d6 2.d4 Nf6 3.Nc3 g6 4.f4
B09.2=Pirc: �sterrikisk attack, 4.f4 Bg7
B09.3=Pirc: �sterrikisk, Ljubojevicvarianten
B09.4=Pirc: �sterrikisk, 5.Nf3
B09.5=Pirc: �sterrikisk, 5...O-O
B09.6=Pirc: �sterrikisk, 5...O-O 6.e5
B09.7=Pirc: �sterrikisk, 5...O-O 6.Be3
B09.8=Pirc: �sterrikisk, 5...O-O 6.Be2
B09.9=Pirc: �sterrikisk, 5...O-O 6.Bd3
B09.10=Pirc: �sterrikisk, 5...O-O 6.Bd3 Nc6
B09.11=Pirc: �sterrikisk, 5...O-O 6.Bd3 Nc6 7.e5
B09.12=Pirc: �sterrikisk, 5...O-O 6.Bd3 Na6
B09.13=Pirc: �sterrikisk, 5...O-O 6.Bd3 Na6 7.O-O c5
B09.14=Pirc: �sterrikisk, 5...O-O 6.Bd3 Na6 7.O-O c5 8.d5
B09.15=Pirc: �sterrikisk, 5...O-O 6.Bd3 Na6 7.O-O c5 8.d5 Bg4
B09.16=Pirc: �sterrikisk, 5...c5
B09.17=Pirc: �sterrikisk, 5...c5 6.dxc5
B09.18=Pirc: �sterrikisk, 5...c5 6.dxc5 Qa5 7.Bd3
B09.19=Pirc: �sterrikisk, 5...c5 6.Bb5+
B09.20=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7
B09.21=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7 7.e5
B09.22=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7 7.e5 Ng4
B09.23=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7 7.e5 Ng4 8.Bxd7+
B09.24=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7 7.e5 Ng4 8.e6
B09.25=Pirc: �sterrikisk, 5...c5, Seirawanvarianten
B09.26=Pirc: �sterrikisk, 5...c5 6.Bb5+ Bd7 7.e5 Ng4 8.e6 Bxb5
B10.1=Caro-Kann: 1.e4 c6
B10.2=Caro-Kann: 2.Ne2
B10.3=Caro-Kann: 2.f4
B10.4=Caro-Kann: Breyervarianten, 1.e4 c6 2.d3
B10.5=Caro-Kann: Breyer, 3.Nd2 g6
B10.6=Caro-Kann: Breyer, 3.Nd2 e5
B10.7=Caro-Kann: Breyer, Huvudvarianten
B10.8=Caro-Kann: Engelska varianten, 2.c4
B10.9=Caro-Kann: Engelska varianten, 2.c4 e5
B10.10=Caro-Kann: Engelska varianten, 2.c4 d5
B10.11=Caro-Kann: Engelska varianten, 2.c4 d5 3.cxd5
B10.12=Caro-Kann: Engelska varianten, 2.c4 d5 3.cxd5 cxd5
B10.13=Caro-Kann: Engelska varianten, 2.c4 d5 3.exd5
B10.14=Caro-Kann: Engelska varianten, 2.c4 d5 3.exd5 cxd5
B10.15=Caro-Kann: Engelskt, Avbyte, 1.e4 c6 2.c4 d5 3.exd5 cxd5 4.cxd5
B10.16=Caro-Kann: Engelskt, Avbyte, 4...Nf6
B10.17=Caro-Kann: Engelskt, Avbyte, 4...Nf6 5.Bb5+
B10.18=Caro-Kann: Engelskt, Avbyte, 4...Nf6 5.Nc3
B10.19=Caro-Kann: 2.Nf3
B10.20=Caro-Kann: 2.Nc3
B10.21=Caro-Kann: 2.Nc3 d5
B10.22=Caro-Kann: Goldman-Spielmann
B10.23=Caro-Kann: Tv� springare-varianten
B10.24=Caro-Kann: Tv� springare, 3...dxe4
B10.25=Caro-Kann: Hectors gambit
B10.26=Caro-Kann: Tv� springare, 3...dxe4 4.Nxe4
B10.27=Caro-Kann: Tv� springare, 3...dxe4 4.Nxe4 Nf6
B11.1=Caro-Kann: Tv� springare, 3...Bg4
B11.2=Caro-Kann: Tv� springare, 3...Bg4 4.h3
B11.3=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bh5
B11.4=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bh5, 7.g4 Bg6
B11.5=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3
B11.6=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3
B11.7=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 dxe4
B11.8=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 dxe4 6.Nxe4
B11.9=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 Nf6
B11.10=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6
B11.11=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d4
B11.12=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.g3
B11.13=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.g3 Nf6
B11.14=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d3
B11.15=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d3 Nd7
B11.16=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d3 Nf6
B11.17=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d3 Nf6 7.a3
B11.18=Caro-Kann: Tv� springare, 3...Bg4 4.h3 Bxf3 5.Qxf3 e6 6.d3 Nf6 7.Bd2
B12.1=Caro-Kann: 2.d4
B12.2=Caro-Kann: de Bruyckers f�rsvar, 1.e4 c6 2.d4 Na6
B12.3=Caro-Kann: Masis f�rsvar, 1.e4 c6 2.d4 Nf6
B12.4=Caro-Kann: 2.d4 d5
B12.5=Caro-Kann: Ulysses gambit, 1.e4 c6 2.d4 d5 3.Nf3
B12.6=Caro-Kann: Ulysses gambit, 3.Nf3 dxe4 4.Ng5
B12.7=Caro-Kann: Mieses gambit, 1.e4 c6 2.d4 d5 3.Be3
B12.8=Caro-Kann: Maroczys (Fantasy)varianten
B12.9=Caro-Kann: Maroczys (Fantasy)varianten, 3...e6
B12.10=Caro-Kann: Maroczys (Fantasy)varianten, 3...dxe4
B12.11=Caro-Kann: Maroczys (Fantasy)varianten, gambitvarianten
B12.12=Caro-Kann: 3.Nd2
B12.13=Caro-Kann: 3.Nd2 dxe4
B12.14=Caro-Kann: Edinburghvarianten, 1.e4 c6 2.d4 d5 3.Nd2 Qb6
B12.15=Caro-Kann: Gurgenidze-Modern: 3.Nd2 g6
B12.16=Caro-Kann: Gurgenidze-Modern: 3.Nd2 g6 4.Ngf3
B12.17=Caro-Kann: Gurgenidze-Modern: 3.Nd2 g6 4.Ngf3 Bg7
B12.18=Caro-Kann: Gurgenidze-Modern: 3.Nd2 g6 4.Ngf3 Bg7 5.h3
B12.19=Caro-Kann: Gurgenidze-Modern: 3.Nd2 g6 4.Ngf3 Bg7 5.c3
B12.20=Caro-Kann: Avanceravarianten, 1.e4 c6 2.d4 d5 3.
B12.21=Caro-Kann: Avanceravarianten, 3...c5
B12.22=Caro-Kann: Avanceravarianten, 3...c5 4.dxc5
B12.23=Caro-Kann: Avanceravarianten, 3...c5 4.dxc5 Nc6
B12.24=Caro-Kann: Avancera, 3...Bf5
B12.25=Caro-Kann: Avancera, Barjonettvarianten
B12.26=Caro-Kann: Avancera, 4.h4
B12.27=Caro-Kann: Avancera, 4.c3
B12.28=Caro-Kann: Avancera, Shortvarianten
B12.29=Caro-Kann: Avancera, 4.Bd3
B12.30=Caro-Kann: Avancera, 4.Nf3
B12.31=Caro-Kann: Avancera, 4.Nf3 e6
B12.32=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2
B12.33=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 Nd7
B12.34=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5
B12.35=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.O-O
B12.36=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.O-O Ne7
B12.37=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.O-O Nd7
B12.38=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.Be3
B12.39=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.Be3 Ne7
B12.40=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.Be3 Nd7
B12.41=Caro-Kann: Avancera, 4.Nf3 e6 5.Be2 c5 6.Be3 Nd7 7.O-O
B12.42=Caro-Kann: Avancera, 4.Nc3
B12.43=Caro-Kann: Avancera, 4.Nc3 h5
B12.44=Caro-Kann: Avancera, 4.Nc3 Qb6
B12.45=Caro-Kann: Avancera, 4.Nc3 e6
B12.46=Caro-Kann: Avancera, Huvudvarianten, 1.e4 c6 2.d4 d5 3.e5 Bf5 4.Nc3 e6 5.g4
B12.47=Caro-Kann: Avancera, Huvudvarianten, 6.Nge2
B12.48=Caro-Kann: Avancera, Huvudvarianten, 6.Nge2 c5
B13.1=Caro-Kann: Avbytesvarianten, 1.e4 c6 2.d4 d5 3.exd5
B13.2=Caro-Kann: Avbyte, 3...Qxd5
B13.3=Caro-Kann: Avbyte, 3...cxd5
B13.4=Caro-Kann: Avbyte, 4.Nf3
B13.5=Caro-Kann: Avbyte, 4.Nf3 Nf6
B13.6=Caro-Kann: Avbyte, 4.Bd3
B13.7=Caro-Kann: Avbyte, 4.Bd3 Nc6
B13.8=Caro-Kann: Avbyte, 4.Bd3 Nc6 5.c3
B13.9=Caro-Kann: Avbyte, 4.Bd3 Nc6 5.c3 g6
B13.10=Caro-Kann: Avbyte, 4.Bd3 Nc6 5.c3 Nf6
B13.11=Caro-Kann: Avbyte, 4.Bd3 Nc6 5.c3 Nf6 6.Nf3
B13.12=Caro-Kann: Avbyte, Rubinsteinvarianten
B13.13=Caro-Kann: Avbyte, Rubinstein, 6...Bg4
B13.14=Caro-Kann: Avbyte, Rubinstein, 7.Qb3 Qc8
B13.15=Caro-Kann: Avbyte, Rubinstein, 7.Qb3 Qd7
B13.16=Caro-Kann: Panov-Botvinnik attack
B13.17=Caro-Kann: Panov-Botvinnik, 4...e6
B13.18=Caro-Kann: Panov-Botvinnik, 4...Nf6
B13.19=Caro-Kann: Panov-Botvinnik, Gunderamvarianten
B13.20=Caro-Kann: Panov-Botvinnik, 5.Nc3
B13.21=Caro-Kann: Panov-Botvinnik, 5...dxc4
B13.22=Caro-Kann: Panov-Botvinnik, 5...dxc4 6.Bxc4
B13.23=Caro-Kann: Panov-Botvinnik, 5...Nc6
B13.24=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.cxd5
B13.25=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.cxd5 Nxd5
B13.26=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3
B13.27=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3 Bg4
B13.28=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3 Bg4 7.cxd5
B13.29=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3 Bg4 7.cxd5 Nxd5
B13.30=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3 Bg4 7.cxd5 Nxd5 8.Qb3
B13.31=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Nf3 Bg4 7.cxd5 Nxd5 8.Qb3 Bxf3 9.gxf3 Nb6
B13.32=Caro-Kann: Panov-Botvinnik, Huvudvarianten, 5...Nc6 6.Nf3 Bg4 7.cxd5 Nxd5 8.Qb3 Bxf3 9.gxf3 e6
B13.33=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Bg5
B13.34=Caro-Kann: Panov-Botvinnik, 5...Nc6, Spielmannarianten
B13.35=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Bg5 dxc4
B13.36=Caro-Kann: Panov-Botvinnik, 5...Nc6, Herzogs f�rsvar
B13.37=Caro-Kann: Panov-Botvinnik, 5...Nc6, Czerniakvarianten
B13.38=Caro-Kann: Panov-Botvinnik, 5...Nc6 6.Bg5 Be6
B13.39=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 1.e4 c6 2.d4 d5 3.exd5 cxd5 4.c4 Nf6 5.Nc3 Nc6 6.Bg5 e6
B13.40=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 7.Nf3
B13.41=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 7.Nf3 Be7
B13.42=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 7.Nf3 Be7 8.c5
B13.43=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 7.Nf3 Be7 8.c5 O-O
B13.44=Caro-Kann: Panov-Botvinnik, 5...Nc6, Normalvarianten, 7.Nf3 Be7 8.c5 O-O 9.Bb5
B14.1=Caro-Kann: Panov-Botvinnik, 5...g6
B14.2=Caro-Kann: Panov-Botvinnik, 5...g6 6.Nf3
B14.3=Caro-Kann: Panov-Botvinnik, 5...g6 6.cxd5
B14.4=Caro-Kann: Panov-Botvinnik, 5...g6 6.cxd5 Nxd5
B14.5=Caro-Kann: Panov-Botvinnik, 5...g6 6.cxd5 Nxd5 7.Bc4
B14.6=Caro-Kann: Panov-Botvinnik, 5...g6 6.cxd5 Bg7
B14.7=Caro-Kann: Panov-Botvinnik, 5...g6 6.Qb3
B14.8=Caro-Kann: Panov-Botvinnik, 5...g6 6.Qb3 Bg7 7.cxd5
B14.9=Caro-Kann: Panov-Botvinnik, 5...g6, Huvudvarianten
B14.10=Caro-Kann: Panov-Botvinnik, 5...g6, Huvudvarianten, 8.Be2
B14.11=Caro-Kann: Panov-Botvinnik, 5...g6, Huvudvarianten, 8.Be2 Nbd7
B14.12=Caro-Kann: Panov-Botvinnik, 5...e6
B14.13=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3
B14.14=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Nc6
B14.15=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Be7
B14.16=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Be7 7.Bd3
B14.17=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Be7 7.cxd5
B14.20=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4
B14.21=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 exd5
B14.22=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5
B14.23=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Qc2
B14.24=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Qc2 Nc6
B14.25=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Qc2 Nc6 9.Bd3
B14.26=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Bd2
B14.27=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Bd2 Nc6
B14.28=Caro-Kann: Panov-Botvinnik, 5...e6 6.Nf3 Bb4 7.cxd5 Nxd5 8.Bd2 Nc6 9.Bd3 O-O
B15.1=Caro-Kann:  1.e4 c6 2.d4 d5 3.Nc3
B15.2=Caro-Kann: Gurgenidze motattack
B15.3=Caro-Kann: Gurgenidze-Modern
B15.4=Caro-Kann: Gurgenidze: 4.Be3
B15.5=Caro-Kann: Gurgenidze: 4.Be3 Bg7
B15.6=Caro-Kann: Gurgenidze: 4.h3
B15.7=Caro-Kann: Gurgenidze: 4.h3 Bg7
B15.8=Caro-Kann: Gurgenidze: 4.e5
B15.9=Caro-Kann: Gurgenidze: 4.e5 Bg7
B15.10=Caro-Kann: Gurgenidze: 4.e5 Bg7 5.f4
B15.11=Caro-Kann: Gurgenidze: 4.e5 Bg7 5.f4 Nh6
B15.12=Caro-Kann: Gurgenidze: 4.e5 Bg7 5.f4 h5
B15.13=Caro-Kann: Gurgenidze: 4.e5 Bg7 5.f4 h5 6.Nf3
B15.14=Caro-Kann: Gurgenidze: 4.Nf3
B15.15=Caro-Kann: Gurgenidze: 4.Nf3 Bg7
B15.16=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.exd5
B15.17=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.e5
B15.18=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.h3
B15.19=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.h3 dxe4
B15.20=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.h3 dxe4 6.Nxe4
B15.21=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.h3 Nf6
B15.22=Caro-Kann: Gurgenidze: 4.Nf3 Bg7 5.h3 Nf6 6.e5
B15.23=Caro-Kann: 3.Nc3 dxe4
B15.24=Caro-Kann: Rasa-Studiers gambit
B15.25=Caro-Kann: von Hennigs gambit
B15.26=Caro-Kann: 4.Nxe4
B15.27=Caro-Kann: 4.Nxe4 Nf6
B15.28=Caro-Kann: 4.Nxe4 Nf6 5.f3 gambit
B15.29=Caro-Kann: Alekhines gambit
B15.30=Caro-Kann: 4.Nxe4 Nf6 5.Ng3
B15.31=Caro-Kann: 4.Nxe4 Nf6 5.Nxf6+
B15.32=Caro-Kann: Tartakower (Nimzowitsch)varianten
B15.33=Caro-Kann: Tartakower, Forgacsvarianten
B15.34=Caro-Kann: Tartakower, 6.c3
B16.1=Caro-Kann: Bronstein-Larsen
B16.2=Caro-Kann: Bronstein-Larsen, 6.Qd3
B16.3=Caro-Kann: Bronstein-Larsen, 6.Ne2
B16.4=Caro-Kann: Bronstein-Larsen, 6.Bc4
B16.5=Caro-Kann: Bronstein-Larsen, 6.Nf3
B16.6=Caro-Kann: Bronstein-Larsen, 6.Nf3 Bf5
B16.7=Caro-Kann: Bronstein-Larsen, 6.Nf3 Bg4
B16.8=Caro-Kann: Bronstein-Larsen, 6.Nf3 Bg4 7.Be2 e6
B16.9=Caro-Kann: Bronstein-Larsen, 6.c3
B16.10=Caro-Kann: Bronstein-Larsen, 6.c3 Bf5
B16.11=Caro-Kann: Bronstein-Larsen, 6.c3 Bf5 7.Ne2
B16.12=Caro-Kann: Bronstein-Larsen, 6.c3 Bf5 7.Nf3
B16.13=Caro-Kann: Bronstein-Larsen, 6.c3 Bf5 7.Nf3 Qc7
B16.14=Caro-Kann: Bronstein-Larsen, 6.c3 Bf5 7.Nf3 e6
B17.1=Caro-Kann: Steinitzvarianten
B17.2=Caro-Kann: Steinitz, 5.Nf3
B17.3=Caro-Kann: Steinitz, 5.Nf3 Ngf6
B17.4=Caro-Kann: Steinitz, 5.Nf3 Ngf6 6.Nxf6+
B17.5=Caro-Kann: Steinitz, 5.Nf3 Ngf6 6.Nxf6+ Nxf6 7.Bc4
B17.6=Caro-Kann: Steinitz, 5.Nf3 Ngf6 6.Ng3
B17.7=Caro-Kann: Steinitz, 5.Nf3 Ngf6 6.Ng3 e6
B17.8=Caro-Kann: Steinitz, 5.Ng5
B17.9=Caro-Kann: Steinitz, 5.Ng5 Ngf6
B17.10=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3
B17.11=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3 e6
B17.12=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3 e6 7.N1f3 Bd6 8.Qe2
B17.13=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3, Huvudvarianten 10.Qxe4
B17.14=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3, Huvudvarianten 10.Qxe4 Qc7
B17.15=Caro-Kann: Steinitz, 5.Ng5 Ngf6 6.Bd3, Huvudvarianten 10.Qxe4 Nf6
B17.16=Caro-Kann: Steinitz, 5.Bc4
B17.17=Caro-Kann: Steinitz, 5.Bc4 Ngf6
B17.18=Caro-Kann: Steinitz, 5.Bc4 Ngf6 6.Ng5
B17.19=Caro-Kann: Steinitz, 5.Bc4 Ngf6 6.Ng5, 8.Bb3
B17.20=Caro-Kann: Steinitz, 5.Bc4 Ngf6 6.Ng5, 8.Bd3
B17.21=Caro-Kann: Steinitz, 5.Bc4 Ngf6 6.Ng5, 8.Bd3 h6
B18.1=Caro-Kann: Klassisk, 1.e4 c6 2.d4 d5 3.Nc3 dxe4 4.Nxe4 Bf5
B18.2=Caro-Kann: Klassisk, 5.Nc5
B18.3=Caro-Kann: Klassisk, 5.Nc5 b6
B18.4=Caro-Kann: Klassisk, 5.Ng3
B18.5=Caro-Kann: Klassisk, 5.Ng3 Bg6
B18.6=Caro-Kann: Klassisk, Maroczy attack
B18.7=Caro-Kann: Klassisk, Flohrvarianten
B18.8=Caro-Kann: Klassisk, 6.N1e2
B18.9=Caro-Kann: Klassisk, 6.Bc4
B18.10=Caro-Kann: Klassisk, 6.Bc4 e6 7.N1e2
B18.11=Caro-Kann: Klassisk, 6.Bc4 e6 7.N1e2 Nf6
B18.12=Caro-Kann: Klassisk, 6.Nf3
B18.13=Caro-Kann: Klassisk, 6.Nf3 Nd7
B18.14=Caro-Kann: Klassisk, 6.Nf3 Nd7 7.Bd3
B18.15=Caro-Kann: Klassisk, 6.Nf3 Nd7 7.Bd3 e6
B18.16=Caro-Kann: Klassisk, 6.h4
B18.17=Caro-Kann: Klassisk, 6.h4 h6
B18.18=Caro-Kann: Klassisk, 6.h4 h6 7.Nh3
B18.19=Caro-Kann: Klassisk, 6.h4 h6 7.f4
B18.20=Caro-Kann: Klassisk, 6.h4 h6 7.h5
B19.1=Caro-Kann: Klassisk, 7.Nf3
B19.2=Caro-Kann: Klassisk, 7.Nf3 e6
B19.3=Caro-Kann: Klassisk, 7.Nf3 Nf6
B19.4=Caro-Kann: Klassisk, 7.Nf3 Nf6 8.h5
B19.5=Caro-Kann: Klassisk, 7.Nf3 Nf6 8.h5
B19.6=Caro-Kann: Klassisk, 7.Nf3 Nf6 8.Ne5
B19.7=Caro-Kann: Klassisk, 7.Nf3 Nf6 8.Ne5 Bh7 9.Bd3
B19.8=Caro-Kann: Klassisk, 7.Nf3 Nd7
B19.9=Caro-Kann: Klassisk, Spasskyvarianten
B19.10=Caro-Kann: Klassisk, Spasskyvarianten
B19.11=Caro-Kann: Klassisk, Spassky, 10.Qxd3
B19.12=Caro-Kann: Klassisk, Spassky, 10.Qxd3 Ngf6
B19.13=Caro-Kann: Klassisk, Spassky, 10.Qxd3 e6
B19.14=Caro-Kann: Klassisk, Spassky, 10.Qxd3 e6 11.Bf4
B19.15=Caro-Kann: Klassisk, Spassky, 10.Qxd3 Qc7
B19.16=Caro-Kann: Klassisk, Spassky, 10.Qxd3 Qc7 11.Bd2
B19.17=Caro-Kann: Klassisk, Spassky, 10.Qxd3 Qc7 11.Bd2 e6
B19.18=Caro-Kann: Klassisk, Spassky, 10.Qxd3 Qc7 11.Bd2 e6 12.O-O-O
B19.19=Caro-Kann: Klassisk, Spassky, Huvudvarianten
B19.20=Caro-Kann: Klassisk, Spassky, Huvudvarianten, 13.Ne4
B19.21=Caro-Kann: Klassisk, Spassky, Huvudvarianten, 13.Ne4 O-O-O
B19.22=Caro-Kann: Klassisk, Spassky, Huvudvarianten, 14.g3 Nxe4
B20.1=Sicilianskt f�rsvar: 1.e4 c5
B20.2=Sicilianskt: Mengarini: 1.e4 c5 2.a3
B20.3=Sicilianskt: Keresvarianten (2.Ne2)
B20.4=Sicilianskt: 2.Bc4
B20.5=Sicilianskt: Vinggambit, 1.e4 c5 2.b4
B20.6=Sicilianskt: Vinggambit, Santasierevarianten, 1.e4 c5 2.b4 cxb4 3.c4
B20.7=Sicilianskt: Vinggambit, Marshallvarianten, 1.e4 c5 2.b4 cxb4 3.a3
B20.8=Sicilianskt: Vinggambit, Marienbadvarianten, 1.e4 c5 2.b4 cxb4 3.a3 d5 4.exd5 Qxd5 5.Bb2
B20.9=Sicilianskt: Vinggambit, Carlsbadvarianten, 1.e4 c5 2.b4 cxb4 3.a3 bxa3
B20.10=Sicilianskt: Snyder, 1.e4 c5 2.b3
B20.11=Sicilianskt: Snyder, 2...e6
B20.12=Sicilianskt: Snyder, 2...d6
B20.13=Sicilianskt: Snyder, 2...Nc6
B20.14=Sicilianskt: Engelskt (2.c4)
B20.15=Sicilianskt: Engelskt, 2...e6
B20.16=Sicilianskt: Engelskt, 2...d6
B20.17=Sicilianskt: Engelskt, 2...Nc6
B20.18=Sicilianskt: Engelskt, 2...Nc6 3.Nf3
B20.19=Sicilianskt: Engelskt, 2...Nc6 3.Ne2
B20.20=Sicilianskt: Engelskt, 2...Nc6 3.Nc3
B20.21=Sicilianskt: Engelskt, 2...Nc6 3.Nc3 g6
B20.22=Sicilianskt: 2.g3
B20.23=Sicilianskt: 2.g3 g6
B20.24=Sicilianskt: 2.g3 g6 3.Bg2 Bg7
B20.25=Sicilianskt: 2.g3 g6 3.Bg2 Bg7 4.f4
B20.26=Sicilianskt: 2.g3 g6 3.Bg2 Bg7 4.f4 d6
B20.27=Sicilianskt: 2.d3
B20.28=Sicilianskt: 2.d3 e6
B20.29=Sicilianskt: 2.d3 e6 3.g3
B20.30=Sicilianskt: 2.d3 Nc6
B20.31=Sicilianskt: 2.d3 Nc6 3.g3
B21.1=Sicilianskt: Grand Prix attack
B21.2=Sicilianskt: Grand Prix, 2...g6
B21.3=Sicilianskt: Grand Prix, 2...d6
B21.4=Sicilianskt: Grand Prix, 2...e6
B21.5=Sicilianskt: Grand Prix, 2...e6 3.Nf3
B21.6=Sicilianskt: Grand Prix, 2...Nc6
B21.7=Sicilianskt: Grand Prix, 2...Nc6 3.d3
B21.8=Sicilianskt: Grand Prix, 2...Nc6 3.Nf3
B21.9=Sicilianskt: Grand Prix, 2...Nc6 3.Nf3 e6
B21.10=Sicilianskt: Grand Prix, 2...Nc6 3.Nf3 g6
B21.11=Sicilianskt: Grand Prix, Tals f�rsvar, 1.e4 c5 2.f4 d5
B21.12=Sicilianskt: Grand Prix, Tals f�rsvar, 3.e5
B21.13=Sicilianskt: Grand Prix, Toiletvarianten, 1.e4 c5 2.f4 d5 3.Nc3
B21.14=Sicilianskt: Grand Prix, Tals f�rsvar, 3.exd5
B21.15=Sicilianskt: Grand Prix, Tals f�rsvar, 1.e4 c5 2.f4 d5 3.exd5 Nf6, 3.exd5 Qxd5
B21.16=Sicilianskt: Grand Prix, Tals gambit
B21.17=Sicilianskt: Grand Prix, Tals gambit, 4.Bb5+
B21.18=Sicilianskt: Smith-Morras gambit, 1.e4 c5 2.d4
B21.19=Sicilianskt: Smith-Morra, 1.e4 c5 2.d4 d5
B21.20=Sicilianskt: Smith-Morra, 1.e4 c5 2.d4 cxd4
B21.21=Sicilianskt: Halasz gambit, 1.e4 c5 2.d4 cxd4 3.f4
B21.22=Sicilianskt: Smith-Morra, Morphy gambit, 1.e4 c5 2.d4 cxd4 3.Nf3
B21.23=Sicilianskt: Smith-Morra, Andreaschek gambit
B21.24=Sicilianskt: Smith-Morra, 3.c3
B21.25=Sicilianskt: Smith-Morra, 3.c3 Nf6
B21.26=Sicilianskt: Smith-Morra, 3.c3 d5
B21.27=Sicilianskt: Smith-Morra, 3.c3 d3
B21.28=Sicilianskt: Antagen Smith-Morra, 1.e4 c5 2.d4 cxd4 3.c3 dxc3
B21.29=Sicilianskt: Antagen Smith-Morra, 1.e4 c5 2.d4 cxd4 3.c3 dxc3 4.Nxc3
B21.30=Sicilianskt: Smith-Morra, 4.Nxc3 d6
B21.31=Sicilianskt: Smith-Morra, 4.Nxc3 e6
B21.32=Sicilianskt: Smith-Morra, 4.Nxc3 e6 5.Nf3
B21.33=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6
B21.34=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6 5.Nf3
B21.35=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6 5.Nf3 e6
B21.36=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6 5.Nf3 e6 6.Bc4
B21.37=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6 5.Nf3 e6 6.Bc4 a6
B21.38=Sicilianskt: Smith-Morra, 4.Nxc3 Nc6 5.Nf3 d6
B21.39=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4
B21.40=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4 a6
B21.41=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4 e6
B21.42=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4 e6 7.O-O
B21.43=Sicilianskt: Smith-Morra gambit, Chicago f�rsvar
B21.44=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4 e6 7.O-O Nf6
B21.45=Sicilianskt: Smith-Morra, 5.Nf3 d6 6.Bc4 e6 7.O-O Nf6 8.Qe2 Be7
B22.1=Sicilianskt: Alapin, 1.e4 c5 2.c3
B22.2=Sicilianskt: Alapin, 2...e5
B22.3=Sicilianskt: Alapin, 2...g6
B22.4=Sicilianskt: Alapin, 2...g6 3.d4
B22.5=Sicilianskt: Alapin, 2...g6 3.d4 cxd4
B22.6=Sicilianskt: Alapin, 2...Nc6
B22.7=Sicilianskt: Alapin, 2...Nc6 3.Nf3
B22.8=Sicilianskt: Alapin, 2...Nc6 3.d4
B22.9=Sicilianskt: Alapin, 2...e6
B22.10=Sicilianskt: Alapin, 2...e6 3.Nf3
B22.12=Sicilianskt: Alapin, 2...e6 3.d4
B22.13=Sicilianskt: Alapin, 2...e6 3.d4 d5
B22.14=Sicilianskt: Alapin, 2...e6 3.d4 d5 4.exd5
B22.15=Sicilianskt: Alapin, 2...e6 3.d4 d5 4.exd5 exd5
B22.16=Sicilianskt: Alapin, 2...e6 3.d4 d5 4.exd5 exd5 5.Nf3
B22.17=Sicilianskt: Alapin, 2...e6 3.d4 d5 4.exd5 exd5 5.Nf3 Nc6
B22.18=Sicilianskt: Alapin, 2...d6
B22.19=Sicilianskt: Alapin, 2...d5
B22.20=Sicilianskt: Alapin, 2...d5 3.exd5
B22.21=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5
B22.22=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4
B22.23=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 cxd4
B22.24=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 cxd4 5.cxd4
B22.25=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 e6
B22.26=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 e6 5.Nf3
B22.27=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nc6
B22.28=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nc6 5.Nf3
B22.29=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nc6 5.Nf3 cxd4
B22.30=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nc6 5.Nf3 cxd4 6.cxd4
B22.31=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nc6 5.Nf3 Bg4
B22.32=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6
B22.33=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6 5.Nf3
B22.34=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6 5.Nf3 Bg4
B22.35=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6 5.Nf3 Bg4 6.Be2 e6
B22.36=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6 5.Nf3 e6 6.Be3
B22.37=Sicilianskt: Alapin, 2...d5 3.exd5 Qxd5 4.d4 Nf6 5.Nf3 e6 6.Be2
B22.38=Sicilianskt: Alapin, 2...Nf6
B22.39=Sicilianskt: Alapin, 2...Nf6 3.e5
B22.40=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5
B22.41=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.g3
B22.42=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.Nf3
B22.43=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.Nf3 Nc6
B22.44=Sicilianskt: Alapin, Heidenfeldvarianten, 1.e4 c5 2.c3 Nf6 3.e5 Nd5 4.Nf3 Nc6 5.Na3
B22.45=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4
B22.46=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4 cxd4
B22.47=Sicilianskt: Alapin, 2...Nf6, 5.Bc4
B22.48=Sicilianskt: Alapin, 2...Nf6, 5.Qxd4
B22.49=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4 cxd4 5.Nf3
B22.50=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4 cxd4 5.Nf3 e6
B22.51=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4 cxd4 5.Nf3 Nc6
B22.52=Sicilianskt: Alapin, 2...Nf6 3.e5 Nd5 4.d4 cxd4 5.Nf3 Nc6 6.Bc4
B22.53=Sicilianskt: Alapin, 2...Nf6, 5.cxd4
B22.54=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 d6
B22.55=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 Nc6
B22.56=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 Nc6 6.Nf3
B22.57=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 d6
B22.58=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 d6 6.Nf3 Nc6
B22.59=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 e6
B22.60=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 e6 6.Nf3
B22.61=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 e6 6.Nf3 Nc6
B22.62=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 e6 6.Nf3 d6
B22.63=Sicilianskt: Alapin, 2...Nf6, 5.cxd4 e6 6.Nf3 b6
B23.1=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3
B23.2=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 g6
B23.3=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 d6
B23.4=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 d6 3.Nge2
B23.5=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 d6 3.g3
B23.6=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 d6 3.f4
B23.7=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 e6
B23.8=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 e6 3.f4
B23.9=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 e6 3.Nge2
B23.10=Sicilianskt: St�ngt, 1.e4 c5 2.Nc3 e6 3.g3
B23.11=Sicilianskt: St�ngt, Korchnoivarianten
B23.12=Sicilianskt: St�ngt, 2...Nc6
B23.13=Sicilianskt: St�ngt, 2...Nc6 3.Bb5
B23.14=Sicilianskt: St�ngt, 2...Nc6 3.Bb5 Nd4
B23.15=Sicilianskt: Chameleonvarianten
B23.16=Sicilianskt: Chameleon, 3...e5
B23.17=Sicilianskt: Chameleon, 3...g6
B23.18=Sicilianskt: St�ngt, Grand Prix
B23.19=Sicilianskt: St�ngt, Grand Prix, 3...d6
B23.20=Sicilianskt: St�ngt, Grand Prix, 3...d6 4.Nf3 g6
B23.21=Sicilianskt: St�ngt, Grand Prix, 3...e6
B23.22=Sicilianskt: St�ngt, Grand Prix, 3...e6 4.Nf3
B23.23=Sicilianskt: St�ngt, Grand Prix, 3...e6 4.Nf3 d5
B23.24=Sicilianskt: St�ngt, Grand Prix, 3...g6
B23.25=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bc4
B23.26=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bc4 e6
B23.27=Sicilianskt: St�ngt, Grand Prix, Schofmanvarianten
B23.28=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bb5
B23.29=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bb5 Nd4
B23.30=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bb5 Nd4 6.Bd3
B23.31=Sicilianskt: St�ngt, Grand Prix, 3...g6 4.Nf3 Bg7 5.Bb5 Nd4 6.O-O
B24.1=Sicilianskt: St�ngt, 3.g3
B24.2=Sicilianskt: St�ngt, 3.g3 e6
B24.3=Sicilianskt: St�ngt, 3.g3 g6
B24.4=Sicilianskt: St�ngt, 3.g3 g6 4.d3
B24.5=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2
B24.6=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7
B24.7=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.Nge2
B24.8=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.f4
B24.9=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.d3
B24.10=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.d3 e6
B24.11=Sicilianskt: St�ngt, Smyslovvarianten
B24.12=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.d3 e6 6.f4
B25.1=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.d3 d6
B25.2=Sicilianskt: St�ngt, 3.g3 g6 4.Bg2 Bg7 5.d3 d6 6.Nge2
B25.3=Sicilianskt: St�ngt, Botvinnik
B25.4=Sicilianskt: St�ngt, 3.g3, 5.d3 d6 6.Nge2 e6
B25.5=Sicilianskt: St�ngt, 6.f4
B25.6=Sicilianskt: St�ngt, 6.f4 Rb8
B25.7=Sicilianskt: St�ngt, 6.f4 Nf6
B25.8=Sicilianskt: St�ngt, 6.f4 Nf6 7.Nf3
B25.9=Sicilianskt: St�ngt, 6.f4 e5
B25.10=Sicilianskt: St�ngt, 6.f4 e5 7.Nf3
B25.11=Sicilianskt: St�ngt, 6.f4 e5 7.Nf3 Nge7
B25.12=Sicilianskt: St�ngt, 6.f4 e5 7.Nf3 Nge7 8.O-O
B25.13=Sicilianskt: St�ngt, 6.f4 e6
B25.14=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3
B25.15=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7
B25.16=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O
B25.17=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O
B25.18=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3
B25.19=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3 Rb8
B25.20=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3 b6
B25.21=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3 Nd4
B25.22=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3 Nd4 10.e5
B25.23=Sicilianskt: St�ngt, 6.f4 e6 7.Nf3 Nge7 8.O-O O-O 9.Be3 Nd4 10.e5 Nef5
B26.1=Sicilianskt: St�ngt, 6.Be3
B26.2=Sicilianskt: St�ngt, 6.Be3 Nf6
B26.3=Sicilianskt: St�ngt, 6.Be3 Nf6 7.h3
B26.4=Sicilianskt: St�ngt, 6.Be3 e5
B26.5=Sicilianskt: St�ngt, 6.Be3 e5 7.Qd2
B26.6=Sicilianskt: St�ngt, 6.Be3 Rb8
B26.7=Sicilianskt: St�ngt, 6.Be3 Rb8 7.Qd2
B26.8=Sicilianskt: St�ngt, 6.Be3 Rb8 7.Qd2 b5
B26.9=Sicilianskt: St�ngt, 6.Be3 Rb8 7.Qd2 b5 8.Nge2
B26.10=Sicilianskt: St�ngt, 6.Be3 e6
B26.11=Sicilianskt: St�ngt, 6.Be3 e6 7.Qd2
B26.12=Sicilianskt: St�ngt, 6.Be3 e6 7.Qd2 Qa5
B26.13=Sicilianskt: St�ngt, 6.Be3 e6 7.Qd2 Nd4
B26.14=Sicilianskt: St�ngt, 6.Be3 e6 7.Qd2 Nge7
B26.15=Sicilianskt: St�ngt, 6.Be3 e6 7.Qd2 Rb8
B27.1=Sicilianskt: 1.e4 c52.Nf3
B27.2=Sicilianskt: Mongoosevarianten
B27.3=Sicilianskt: Quinterosvarianten
B27.4=Sicilianskt: Katalimovvarianten
B27.5=Sicilianskt: Ungerska varianten, 1.e4 c5 2.Nf3 g6
B27.6=Sicilianskt: Ungersk, 3.c4
B27.7=Sicilianskt: Ungersk, 3.c3
B27.8=Sicilianskt: Ungersk, 3.c3 Bg7 4.d4 cxd4 5.cxd4
B27.9=Sicilianskt: Ungersk, 3.d4
B27.10=Sicilianskt: Ungersk, 3.d4 cxd4
B27.11=Sicilianskt: Ungersk, 3.d4 cxd4 4.Nxd4
B27.12=Sicilianskt: Accelererad Pterodactyl, 1.e4 c5 2.Nf3 g6 3.d4 Bg7
B27.13=Sicilianskt: Accelererad Pterodactyl, 4.dxc5
B27.14=Sicilianskt: Accelererad Pterodactyl, 4.dxc5 Qa5+
B27.15=Sicilianskt: Accelererad Pterodactyl, 4.dxc5 Qa5+ 5.Nc3
B27.16=Sicilianskt: Accelererad Pterodactyl, 4.dxc5 Qa5+ 5.c3
B27.17=Sicilianskt: Accelererad Pterodactyl, 4.dxc5 Qa5+ 5.c3
B27.19=Sicilianskt: Accelererad Pterodactyl, 4.Nc3
B28.1=Sicilianskt: O'Kellyvarianten, 1.e4 c5 2.Nf3 a6
B28.2=Sicilianskt: O'Kelly, 3.Nc3
B28.3=Sicilianskt: O'Kelly, 3.d4
B28.4=Sicilianskt: O'Kelly, 3.d4 cxd4 4.Nxd4
B28.5=Sicilianskt: O'Kelly, 3.d4 cxd4 4.Nxd4 Nf6
B28.6=Sicilianskt: O'Kelly, 3.c4
B28.7=Sicilianskt: O'Kelly, 3.c4 e6
B28.8=Sicilianskt: O'Kelly, 3.c3
B28.9=Sicilianskt: O'Kelly, 3.c3 d5
B29.1=Sicilianskt: Nimzowitsch, 1.e4 c5 2.Nf3 Nf6
B29.2=Sicilianskt: Nimzowitsch, 3.d3
B29.3=Sicilianskt: Nimzowitsch, 3.Nc3
B29.4=Sicilianskt: Nimzowitsch, 3.Nc3 d5
B29.5=Sicilianskt: Nimzowitsch, 3.e5
B29.6=Sicilianskt: Nimzowitsch, 3.e5 Nd5
B29.7=Sicilianskt: Nimzowitsch, 4.c4
B29.8=Sicilianskt: Nimzowitsch, 4.d4
B29.9=Sicilianskt: Nimzowitsch, 4.Nc3
B29.10=Sicilianskt: Nimzowitsch, 4.Nc3 Nxc3
B29.11=Sicilianskt: Nimzowitsch, 4.Nc3 e6
B29.12=Sicilianskt: Nimzowitsch, 4.Nc3 e6 5.Nxd5
B29.13=Sicilianskt: Nimzowitsch, Rubinsteins motgambit
B29.14=Sicilianskt: Nimzowitsch, Rubinsteins motgambit, 7.dxc5
B30.1=Sicilianskt: 1.e4 c5 2.Nf3 Nc6
B30.2=Sicilianskt: 2...Nc6 3.b3
B30.3=Sicilianskt: 2...Nc6 3.d3
B30.4=Sicilianskt: 2...Nc6 3.d3 Nf6
B30.5=Sicilianskt: 2...Nc6 3.g3
B30.6=Sicilianskt: 2...Nc6 3.g3 e6 4.d3
B30.8=Sicilianskt: 2...Nc6 3.Bc4
B30.9=Sicilianskt: 2...Nc6 3.Nc3
B30.10=Sicilianskt: 2...Nc6 3.Nc3 Nf6
B30.11=Sicilianskt: 2...Nc6 3.Nc3 g6
B30.12=Sicilianskt: 2...Nc6 3.Nc3 e5
B30.13=Sicilianskt: Rossolimo, 1.e4 c5 2.Nf3 Nc6 3.Bb5
B30.14=Sicilianskt: Rossolimo, 3...Qb6
B30.15=Sicilianskt: Rossolimo, 3...Nf6
B30.16=Sicilianskt: Rossolimo, 3...e6
B30.17=Sicilianskt: Rossolimo, 3...e6 4.b3
B30.18=Sicilianskt: Rossolimo, 3...e6 4.Nc3
B30.19=Sicilianskt: Rossolimo, 3...e6 4.Bxc6
B30.20=Sicilianskt: Rossolimo, 3...e6 4.O-O
B30.21=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7
B30.22=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7 5.b3
B30.23=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7 5.Re1
B30.24=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7 5.Nc3
B30.25=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7 5.c3
B30.26=Sicilianskt: Rossolimo, 3...e6 4.O-O Nge7 5.c3 a6
B31.1=Sicilianskt: Rossolimo, 1.e4 c5 2.Nf3 Nc6 3.Bb5 g6
B31.2=Sicilianskt: Rossolimo, 3...g6 4.Nc3
B31.3=Sicilianskt: Rossolimo, 3...g6 4.Bxc6
B31.4=Sicilianskt: Rossolimo, 3...g6 4.Bxc6 dxc6
B31.5=Sicilianskt: Rossolimo, 3...g6 4.Bxc6 dxc6 5.d3
B31.6=Sicilianskt: Rossolimo, 3...g6 4.Bxc6 dxc6 5.d3 Bg7 6.h3
B31.7=Sicilianskt: Rossolimo, 3...g6 4.O-O
B31.8=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.c3
B31.9=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.c3 e5
B31.10=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1
B31.11=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 Nf6
B31.12=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 Nf6 6.c3
B31.13=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 Nf6 6.c3 O-O 7.h3
B31.14=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 Nf6 6.c3 O-O 7.d4
B31.15=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 e5
B31.16=Sicilianskt: Rossolimo, Gurgenidzevarianten
B31.17=Sicilianskt: Rossolimo, 3...g6 4.O-O Bg7 5.Re1 e5
B32.1=Sicilianskt: 1.e4 c5 2.Nf3 Nc6 3.d4
B32.2=Sicilianskt: 2...Nc6 3.d4 cxd4
B32.3=Sicilianskt: �ppet, 2...Nc6
B32.5=Sicilianskt: �ppet, 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 Qb6
B32.6=Sicilianskt: Flohrvarianten
B32.7=Sicilianskt: Flohr, 5.Nb5
B32.8=Sicilianskt: Nimzowitschvarianten, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 d5
B32.9=Sicilianskt: L�wenthal, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 e5
B32.10=Sicilianskt: L�wenthal, 5.Nb5
B32.11=Sicilianskt: L�wenthal, 5...a6
B32.12=Sicilianskt: L�wenthal, Dambyte, 5...a6
B32.13=Sicilianskt: L�wenthal, 5...a6, 6.Nd6+ Bxd6 7.Qxd6 Qf6 8.Qd1
B32.14=Sicilianskt: L�wenthal, Kalashnikov, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 e5 5.Nb5 d6
B32.15=Sicilianskt: L�wenthal, Kalashnikov, 6.a4
B32.16=Sicilianskt: L�wenthal, Kalashnikov, 6.N1c3
B32.17=Sicilianskt: L�wenthal, Kalashnikov, 6.N1c3 a6 7.Na3 b5
B32.18=Sicilianskt: L�wenthal, Kalashnikov, 6.N1c3 a6 7.Na3 b5 8.Nd5 Nge7
B32.19=Sicilianskt: L�wenthal, Kalashnikov, 6.c4
B32.20=Sicilianskt: L�wenthal, Kalashnikov, 6.c4 Be7
B32.21=Sicilianskt: L�wenthal, Kalashnikov, 6.c4 Be7 7.Be2
B32.22=Sicilianskt: L�wenthal, Kalashnikov, 6.c4 Be7 7.N1c3
B32.23=Sicilianskt: L�wenthal, Kalashnikov, Huvudvarianten
B32.24=Sicilianskt: L�wenthal, Kalashnikov, Huvudvarianten, 9.Nc2
B32.25=Sicilianskt: L�wenthal, Kalashnikov, Huvudvarianten, 9.Be2
B33.1=Sicilianskt: �ppet, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 Nf6
B33.2=Sicilianskt: �ppet, 2...Nc6, 5...Qb6
B33.3=Sicilianskt: �ppet, 2...Nc6, 5...Qb6 6.Nb3
B33.4=Sicilianskt: �ppet, 2...Nc6, 5...Qb6 6.Nb3 e6
B33.5=Sicilianskt: �ppet, 2...Nc6, 5...Qb6 6.Nb3 e6 7.Bd3
B33.6=Sicilianskt: Pelikan-Sveshnikov, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e5
B33.7=Sicilianskt: Pelikan-Sveshnikov, 6.Nxc6
B33.8=Sicilianskt: Pelikan-Sveshnikov, 6.Nf5
B33.9=Sicilianskt: Pelikan-Sveshnikov, 6.Nf3
B33.10=Sicilianskt: Pelikan-Sveshnikov, 6.Nb3
B33.11=Sicilianskt: Pelikan-Sveshnikov, 6.Nbd5
B33.12=Sicilianskt: Pelikan, Haberditzvarianten, 6.Ndb5 h6
B33.13=Sicilianskt: Pelikan-Sveshnikov, Pelikanvarianten, 6.Ndb5 d6
B33.14=Sicilianskt: Pelikan, 7.Na3
B33.15=Sicilianskt: Pelikan, 7.a4
B33.16=Sicilianskt: Pelikan, 7.a4
B33.17=Sicilianskt: Pelikan, 7.Nd5
B33.18=Sicilianskt: Pelikan, 7.Bg5
B33.19=Sicilianskt: Pelikan, 7.Bg5 a6
B33.20=Sicilianskt: Pelikan, 7.Bg5 a6 8.Bxf6
B33.21=Sicilianskt: Pelikan, 7.Bg5 a6 8.Na3
B33.22=Sicilianskt: Pelikan, Birdvarianten
B33.23=Sicilianskt: Pelikan, Chelyabinskvariant, 8..b5
B33.24=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5
B33.25=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7
B33.26=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7, 11.c3
B33.27=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7, 11.c3 O-O
B33.28=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7, 11.c3 Bg5
B33.29=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7, 11.c3 O-O 12.Nc2 Bg5
B33.30=Sicilianskt: Pelikan, Chelyabinsk, 9.Nd5 Be7, 11.c3 O-O 12.Nc2 Bg5 13.a4
B33.31=Sicilianskt: Pelikan, Chelyabinsk, 9.Bxf6
B33.32=Sicilianskt: Pelikan, Chelyabinsk, 9.Bxf6 gxf6
B33.33=Sicilianskt: Pelikan, Chelyabinsk, 9.Bxf6 gxf6 10.Nd5
B33.34=Sicilianskt: Pelikan, Chelyabinsk, 9.Bxf6 gxf6 10.Nd5 Bg7
B33.35=Sicilianskt: Pelikan, Chelyabinsk, 9.Bxf6 gxf6 10.Nd5 Bg7 11.Bd3
B33.36=Sicilianskt: Pelikan, Sveshnikovvarianten, 10..f5
B33.37=Sicilianskt: Pelikan, Sveshnikov, 11.c3
B33.38=Sicilianskt: Pelikan, Sveshnikov, 11.c3 Bg7
B33.39=Sicilianskt: Pelikan, Sveshnikov, 11.c3 Bg7 12.exf5 Bxf5
B33.40=Sicilianskt: Pelikan, Sveshnikov, 11.c3 Bg7 12.exf5 Bxf5 13.Nc2 O-O
B33.41=Sicilianskt: Pelikan, Sveshnikov, 11.Bd3
B33.42=Sicilianskt: Pelikan, Sveshnikov, 11.Bd3 Be6
B33.43=Sicilianskt: Pelikan, Sveshnikov, 11.Bd3 Be6 12.O-O
B34.1=Sicilianskt: Accelererad Fianchetto, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 g6
B34.2=Sicilianskt: Accelererad Fianchetto, 5.Bc4
B34.3=Sicilianskt: Accelererad Fianchetto, Avbytesvarianten, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 g6 5.Nxc6
B34.4=Sicilianskt: Accelererad Fianchetto, 5.Be2
B34.5=Sicilianskt: Accelererad Fianchetto, 5.Be3
B34.6=Sicilianskt: Accelererad Fianchetto, Modern variant
B34.7=Sicilianskt: Accelererad Fianchetto, Modern, 5...Nf6
B34.8=Sicilianskt: Accelererad Fianchetto, Modern, 5...Nf6 6.Nxc6
B34.9=Sicilianskt: Accelererad Fianchetto, Modern, 5...Nf6 6.Nxc6 bxc6
B34.10=Sicilianskt: Accelererad Fianchetto, Modern, 5...Bg7
B34.11=Sicilianskt: Accelererad Fianchetto, Modern, 6.Nde2
B34.12=Sicilianskt: Accelererad Fianchetto, Modern, 6.Nb3
B34.13=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3
B34.14=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 d6
B34.15=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 d6 7.Qd2
B34.16=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6
B34.17=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.f3
B34.18=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Nxc6
B34.19=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Nxc6 bxc6
B34.20=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Nxc6 bxc6 8.e5
B34.21=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Nxc6 bxc6 8.e5 Ng8
B34.22=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Be2
B34.23=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Be2 O-O
B34.24=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Be2 O-O 8.O-O
B34.25=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Be2 O-O 8.O-O d5
B34.26=Sicilianskt: Accelererad Fianchetto, Modern, 6.Be3 Nf6 7.Be2 O-O 8.O-O d5 9.exd5
B35.1=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4
B35.2=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 Qa5
B35.3=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 Qa5 8.O-O O-O
B35.4=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 Qa5 8.O-O O-O 9.Bb3
B35.5=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 Qa5 8.O-O O-O 9.Bb3 d6 10.h3 Bd7 11.f4
B35.6=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O
B35.7=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.f3
B35.8=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.O-O
B35.9=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3
B35.10=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3 Ng4
B35.11=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3 Qa5
B35.12=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3 a5
B35.13=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3 a5 9.a4
B35.14=Sicilianskt: Accelererad Fianchetto, Modern, 7.Bc4 O-O 8.Bb3 a5 9.f3
B36.1=Sicilianskt: Maroczy Bind, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 g6 5.c4
B36.2=Sicilianskt: Maroczy Bind, 5...d6
B36.3=Sicilianskt: Maroczy Bind, 5...d6 6.Nc3
B36.4=Sicilianskt: Maroczy Bind, 5...d6 6.Nc3 Bg7
B36.5=Sicilianskt: Maroczy Bind, 5...Nf6
B36.6=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3
B36.7=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 Nxd4
B36.8=Sicilianskt: Maroczy Bind, Gurgenidzevarianten
B36.9=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6
B36.10=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2
B36.11=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4
B36.12=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7
B36.13=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.O-O
B36.14=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Bg5
B36.15=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Bg5 O-O
B36.16=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Bg5 O-O 10.Qd2
B36.17=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Be3
B36.18=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Be3 O-O
B36.19=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Be3 O-O 10.Qd2
B36.20=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Be3 O-O 10.Qd2 Be6
B36.21=Sicilianskt: Maroczy Bind, 5...Nf6 6.Nc3 d6 7.Be2 Nxd4 8.Qxd4 Bg7 9.Be3 O-O 10.Qd2 Be6 11.O-O
B37.1=Sicilianskt: Maroczy Bind, 5...Bg7
B37.2=Sicilianskt: Maroczy Bind, 6.Nb3
B37.3=Sicilianskt: Maroczy Bind, 6.Nc2
B37.4=Sicilianskt: Maroczy Bind, 6.Nc2 d6
B37.5=Sicilianskt: Maroczy Bind, 6.Nc2 d6 7.Be2
B37.6=Sicilianskt: Maroczy Bind, Simaginvarianten
B37.7=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6
B37.8=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3
B37.9=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 O-O
B37.10=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6
B37.11=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2
B37.12=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 Nd7
B37.13=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O
B37.14=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O
B37.15=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Be6
B37.16=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Nd7
B37.17=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Nd7 10.Bd2
B37.18=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Nd7 10.Bd2 a5
B37.19=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Nd7 10.Bd2 Nc5
B37.20=Sicilianskt: Maroczy Bind, 6.Nc2 Nf6 7.Nc3 d6 8.Be2 O-O 9.O-O Nd7 10.Bd2 Nc5 11.b4
B38.1=Sicilianskt: Maroczy Bind, 6.Be3
B38.2=Sicilianskt: Maroczy Bind, 6.Be3 Nh6
B38.3=Sicilianskt: Maroczy Bind, 6.Be3 d6
B38.4=Sicilianskt: Maroczy Bind, 6.Be3 d6 7.Nc3 Nh6
B38.5=Sicilianskt: Maroczy Bind, 6.Be3 Nf6
B38.6=Sicilianskt: Maroczy Bind, 6.Be3 Nf6 7.Nc3
B38.7=Sicilianskt: Maroczy Bind, 6.Be3 Nf6 7.Nc3 d6
B38.8=Sicilianskt: Maroczy Bind, 6.Be3 Nf6 7.Nc3 d6 8.Be2
B38.9=Sicilianskt: Maroczy Bind, 7.Nc3 O-O
B38.10=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2
B38.11=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 b6
B38.12=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 b6 9.O-O
B38.13=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 b6 9.O-O Bb7
B38.14=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 b6 9.O-O Bb7 10.f3
B38.15=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 b6 9.O-O Bb7 10.f3 Qb8
B38.16=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6
B38.17=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.f3
B38.18=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O
B38.19=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Nd7
B38.20=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O a6
B38.21=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Nxd4
B38.22=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7
B38.23=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Nc2
B38.24=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.f3
B38.25=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Rc1
B38.26=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2
B38.27=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2 Nxd4
B38.28=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2 Nxd4 11.Bxd4
B38.29=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2 Nxd4, 12.f3
B38.30=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2 Nxd4, 12.f3 a5
B38.31=Sicilianskt: Maroczy Bind, 7.Nc3 O-O 8.Be2 d6 9.O-O Bd7 10.Qd2 Nxd4, 12.f3 a5 13.b3
B39.1=Sicilianskt: Maroczy Bind, Breyervarianten, 1.e4 c5 2.Nf3 Nc6 3.d4 cxd4 4.Nxd4 g6 5.c4 Bg7 6.Be3 Nf6 7.Nc3 Ng4
B39.2=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4
B39.3=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4
B39.4=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1
B39.5=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 e5
B39.6=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 e5 10.Nb5
B39.7=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 e5 10.Bd3
B39.8=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 Ne6
B39.9=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 Ne6 10.Qd2
B39.10=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 Ne6 10.Rc1
B39.11=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 Ne6 10.Rc1 Qa5
B39.12=Sicilianskt: Maroczy Bind, Breyer, 8.Qxg4 Nxd4 9.Qd1 Ne6 10.Rc1 Qa5 11.Qd2
B40.1=Sicilianskt: 1.e4 c5 2.Nf3 e6
B40.2=Sicilianskt: 2...e6 3.c4
B40.3=Sicilianskt: 2...e6 3.b3
B40.4=Sicilianskt: 2...e6 3.b3 Nc6
B40.5=Sicilianskt: 2...e6 3.g3
B40.6=Sicilianskt: 2...e6 3.d3
B40.7=Sicilianskt: 2...e6 3.Nc3
B40.8=Sicilianskt: 2...e6 3.Nc3 Nc6
B40.9=Sicilianskt: 2...e6 3.d4
B40.10=Sicilianskt: Marshallvarianten, 1.e4 c5 2.Nf3 e6 3.d4 d5
B40.11=Sicilianskt: �ppet, 2...e6
B40.12=Sicilianskt: �ppet, 2...e6, 4.Nxd4
B40.13=Sicilianskt: �ppet, 2...e6, 4.Nxd4 d6
B40.14=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Bc5
B40.15=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Nf6
B40.16=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Nf6 5.Bd3
B40.17=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Nf6 5.Bd3 Nc6
B40.18=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Nf6 5.Bd3 Nc6 6.Nxc6
B40.19=Sicilianskt: �ppet, 2...e6, 4.Nxd4 Nf6 5.Nc3
B40.20=Sicilianskt: Pinvarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Bb4
B40.21=Sicilianskt: Pin, Jaffevarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Bb4 6.Bd3 e5
B40.22=Sicilianskt: Pin, Kochvarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Bb4 6.e5
B41.1=Sicilianskt: Kan (Paulsen) varianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 a6
B41.2=Sicilianskt: Kan, 5.g3
B41.3=Sicilianskt: Kan, 5.Be3
B41.4=Sicilianskt: Kan, 5.Be2
B41.5=Sicilianskt: Kan, 5.Be2 Nf6
B41.6=Sicilianskt: Kan, 5.c4
B41.7=Sicilianskt: Kan, 5.c4 Qc7
B41.8=Sicilianskt: Kan, 5.c4 Nf6
B41.9=Sicilianskt: Kan, 5.c4 Nf6 6.Nc3
B41.10=Sicilianskt: Kan, 5.c4 Nf6 6.Nc3 d6
B41.11=Sicilianskt: Kan, 5.c4 Nf6 6.Nc3 Bb4
B41.12=Sicilianskt: Kan, 5.c4 Nf6, Bronsteinvarianten
B41.13=Sicilianskt: Kan, 5.c4 Nf6 6.Nc3 Qc7
B41.14=Sicilianskt: Kan, 5.c4 Nf6 6.Nc3 Qc7 7.Be2
B42.1=Sicilianskt: Kan, 5.Bd3
B42.2=Sicilianskt: Kan, Schweizisk ostvariant, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 a6 5.Bd3 g6
B42.3=Sicilianskt: Kan, 5.Bd3 Qb6
B42.4=Sicilianskt: Kan, 5.Bd3 Qc7
B42.5=Sicilianskt: Kan, 5.Bd3 Nc6
B42.6=Sicilianskt: Kan, Polugaevskyvarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 a6 5.Bd3 Bc5
B42.7=Sicilianskt: Kan, Polugaevsky, 6.Nb3 Ba7
B42.8=Sicilianskt: Kan, 5.Bd3 Nf6
B42.9=Sicilianskt: Kan, 5.Bd3 Nf6 6.c4
B42.10=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O
B42.11=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O d6
B42.12=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O d6 7.c4
B42.13=Sicilianskt: Kan, Gipslisvarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 a6 5.Bd3 Nf6 6.O-O d6 7.c4 g6
B42.14=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O Qc7
B42.15=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O Qc7 7.c4
B42.16=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O Qc7 7.Qe2
B42.17=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O Qc7 7.Qe2
B42.18=Sicilianskt: Kan, 5.Bd3 Nf6 6.O-O Qc7 7.Qe2 d6 8.c4
B43.1=Sicilianskt: Kan, 5.Nc3
B43.3=Sicilianskt: Kan, 5.Nc3 b5
B43.4=Sicilianskt: Kan, 5.Nc3 b5 6.Bd3
B43.5=Sicilianskt: Kan, 5.Nc3 b5 6.Bd3 Qb6
B43.6=Sicilianskt: Kan, 5.Nc3 b5 6.Bd3 Qb6 7.Nb3
B43.7=Sicilianskt: Kan, 5.Nc3 Qc7
B43.8=Sicilianskt: Kan, 5.Nc3 Qc7 6.g3
B43.9=Sicilianskt: Kan, 5.Nc3 Qc7 6.g3 Nf6
B43.10=Sicilianskt: Kan, 5.Nc3 Qc7 6.Be2
B43.11=Sicilianskt: Kan, 5.Nc3 Qc7 6.Be2 Nf6
B43.12=Sicilianskt: Kan, 5.Nc3 Qc7 6.Be2 Nf6 7.O-O
B43.13=Sicilianskt: Kan, 5.Nc3 Qc7 6.Bd3
B43.14=Sicilianskt: Kan, 5.Nc3 Qc7 6.Bd3 Nf6
B43.15=Sicilianskt: Kan, 5.Nc3 Qc7 6.Bd3 Nf6 7.O-O
B44.1=Sicilianskt: Taimanov, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 Nc6
B44.2=Sicilianskt: Taimanov, 5.g3
B44.3=Sicilianskt: Taimanov, 5.Be2
B44.4=Sicilianskt: Taimanov, 5.c4
B44.5=Sicilianskt: Taimanov, 5.c4 Nf6
B44.6=Sicilianskt: Taimanov, 5.c4 Nf6 6.Nc3
B44.7=Sicilianskt: Taimanov, 5.c4 Nf6 6.Nc3 Bb4
B44.8=Sicilianskt: Taimanov, 5.c4 Nf6 6.Nc3 Bb4 7.Nxc6
B44.9=Sicilianskt: Taimanov, 5.c4 Nf6 6.Nc3 Bb4 7.Nxc6 bxc6
B44.10=Sicilianskt: Taimanov, 5.Be3
B44.11=Sicilianskt: Taimanov, 5.Be3 Nf6
B44.12=Sicilianskt: Taimanov, 5.Nxc6
B44.13=Sicilianskt: Taimanov, 5.Nxc6 bxc6 6.Bd3
B44.14=Sicilianskt, Taimanov, Szenvarianten
B44.15=Sicilianskt, Taimanov, Szen, 5...d6
B44.16=Sicilianskt, Taimanov, Szen, 6.Bf4
B44.17=Sicilianskt, Taimanov, Szen, 6.Bf4 e5 7.Be3 a6
B44.18=Sicilianskt, Taimanov, Szen, 6.Bf4 e5 7.Be3 Nf6
B44.19=Sicilianskt, Taimanov, Szen, 6.c4
B44.20=Sicilianskt, Taimanov, Szen, 6.c4 a6
B44.21=Sicilianskt, Taimanov, Szen, 6.c4 Nf6
B44.22=Sicilianskt, Taimanov, Szen, 7.N5c3
B44.23=Sicilianskt, Taimanov, Szen, 7.N1c3
B44.24=Sicilianskt, Taimanov, Szen, 7.N1c3 a6
B44.25=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3
B44.26=Sicilianskt: Taimanov, Szen, Kasparov gambit, 8.Na3 d5
B44.27=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3 b6
B44.28=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3 Be7
B44.29=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3 Be7 9.Be2
B44.30=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3 Be7 9.Be2 b6
B44.31=Sicilianskt, Taimanov, Szen, 7.N1c3 a6 8.Na3 Be7 9.Be2 O-O
B44.32=Sicilianskt: Taimanov, Szen, Hedgehogvarianten
B44.33=Sicilianskt: Taimanov, Szen, Hedgehog, 11.Be3
B44.34=Sicilianskt: Taimanov, Szen, Hedgehog, 11.Be3 Bd7
B44.35=Sicilianskt: Taimanov, Szen, Hedgehog, 11.Be3 Ne5
B44.36=Sicilianskt: Taimanov, Szen, Hedgehog, 11.Be3 Bb7
B44.37=Sicilianskt: Taimanov, Szen, Hedgehog, 11.Be3 Bb7 12.Qb3
B45.1=Sicilianskt: Taimanov, 5.Nc3
B45.2=Sicilianskt: Taimanov, 5.Nc3 Bb4
B45.5=Sicilianskt: Taimanov, Fyra Springare
B45.6=Sicilianskt: Taimanov, Fyra Springare, 6.Bg5
B45.7=Sicilianskt: Taimanov, Fyra Springare, 6.a3
B45.8=Sicilianskt: Taimanov, Fyra Springare, 6.g3
B45.9=Sicilianskt: Taimanov, Fyra Springare, 6.Be2
B45.10=Sicilianskt: Taimanov, Fyra Springare, 6.Be3
B45.11=Sicilianskt: Taimanov, Fyra Springare, 6.Be3 Bb4
B45.12=Sicilianskt: Taimanov, Fyra Springare, 6.Be3 Bb4 7.Bd3
B45.13=Sicilianskt: Taimanov, Fyra Springare, 6.Nxc6
B45.14=Sicilianskt: Taimanov, Fyra Springare, 6.Nxc6 bxc6 7.e5
B45.15=Sicilianskt: Taimanov, Fyra Springare, 6.Nxc6 bxc6 7.e5 Nd5
B45.16=Sicilianskt: Taimanov, Fyra Springare, 6.Nxc6 bxc6 7.e5 Nd5 8.Ne4
B45.17=Sicilianskt: Taimanov, Fyra Springare, 6.Nxc6 bxc6 7.e5 Nd5 8.Ne4 Qc7
B45.18=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5
B45.19=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 d6
B45.20=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 d6 7.Bf4
B45.21=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4
B45.22=Sicilianskt: Taimanov, Fyra Springare, American attack
B45.23=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3
B45.24=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3 Bxc3+ 8.Nxc3 d5
B45.25=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3, 9.ed5 ed5
B45.26=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3, 9.ed5 ed5 10.Bd3 O-O
B45.27=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3, 10.Bd3 O-O 11.O-O d4
B45.28=Sicilianskt: Taimanov, Fyra Springare, 6.Ndb5 Bb4 7.a3, 10.Bd3 O-O 11.O-O d4 12.Ne2
B46.1=Sicilianskt: Taimanov, 5...a6
B46.2=Sicilianskt: Taimanov, 5...a6 6.f4
B46.3=Sicilianskt: Taimanov, 5...a6 6.Nxc6
B46.4=Sicilianskt: Taimanov, 5...a6 6.Nxc6 bxc6 7.Bd3
B46.5=Sicilianskt: Taimanov, 5...a6 6.Nxc6 bxc6 7.Bd3 d5
B46.6=Sicilianskt: Taimanov, 5...a6 6.g3
B46.7=Sicilianskt: Taimanov, 5...a6 6.g3 Nge7
B46.8=Sicilianskt: Taimanov, 5...a6 6.g3 d6
B46.9=Sicilianskt: Taimanov, 5...a6 6.Be3
B46.10=Sicilianskt: Taimanov, 5...a6 6.Be3 d6
B46.11=Sicilianskt: Taimanov, 5...a6 6.Be3 Nge7
B46.12=Sicilianskt: Taimanov, 5...a6 6.Be3 Nf6
B46.13=Sicilianskt: Taimanov, 5...a6 6.Be2
B46.14=Sicilianskt: Taimanov, 5...a6 6.Be2 Nf6
B46.15=Sicilianskt: Taimanov, 5...a6 6.Be2 Nge7
B46.16=Sicilianskt: Taimanov, 5...a6 6.Be2 Nge7 7.O-O
B46.17=Sicilianskt: Taimanov, 5...a6 6.Be2 Nge7 7.Be3
B47.1=Sicilianskt: Taimanov, Bastrikovvarianten, 1.e4 c5 2.Nf3 e6 3.d4 cxd4 4.Nxd4 Nc6 5.Nc3 Qc7
B47.2=Sicilianskt: Taimanov, 6.Nxc6
B47.3=Sicilianskt: Taimanov, 6.Ndb5
B47.4=Sicilianskt: Taimanov, 6.f4
B47.5=Sicilianskt: Taimanov, 6.f4 a6
B47.6=Sicilianskt: Taimanov, 6.f4 a6 7.Nxc6
B47.7=Sicilianskt: Taimanov, 6.g3
B47.8=Sicilianskt: Taimanov, 6.g3 a6
B47.9=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2
B47.10=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 d6
B47.11=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 d6 8.O-O
B47.12=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 d6 8.O-O Bd7
B47.13=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 d6 8.O-O Bd7 9.Re1
B47.14=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 Nf6
B47.15=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 Nf6 8.O-O
B47.16=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 Nf6 8.O-O Bc5
B47.17=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 Nf6 8.O-O Be7
B47.18=Sicilianskt: Taimanov, 6.g3 a6 7.Bg2 Nf6 8.O-O Be7 9.Re1
B47.19=Sicilianskt: Taimanov, 6.Be2
B47.20=Sicilianskt: Taimanov, 6.Be2 Nf6
B47.21=Sicilianskt: Taimanov, 6.Be2 a6
B47.22=Sicilianskt: Taimanov, 6.Be2 a6 7.f4
B47.23=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O
B47.24=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O b5
B47.25=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6
B47.26=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.a3
B47.27=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1
B47.28=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1 Be7
B47.29=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1 Nxd4
B47.30=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1 Nxd4, 10.Qd3
B47.31=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1 Nxd4, 10.Qd3 b5
B47.32=Sicilianskt: Taimanov, 6.Be2 a6 7.O-O Nf6 8.Kh1 Nxd4, 10.Qd3 b5 11.f4
B48.1=Sicilianskt: Taimanov, 6.Be3
B48.2=Sicilianskt: Taimanov, 6.Be3 Nf6
B48.3=Sicilianskt: Taimanov, 6.Be3 a6
B48.4=Sicilianskt: Taimanov, 6.Be3 a6 7.a3
B48.5=Sicilianskt: Taimanov, 6.Be3 a6 7.f4
B48.6=Sicilianskt: Taimanov, 6.Be3 a6 7.f4 b5
B48.7=Sicilianskt: Taimanov, 6.Be3 a6 7.Qd2
B48.8=Sicilianskt: Taimanov, 6.Be3 a6 7.Qd2 Nf6 8.f3
B48.9=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3
B48.10=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 b5
B48.11=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 b5 8.Nxc6
B48.12=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 b5 8.O-O
B48.13=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6
B48.14=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O
B48.15=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Nxd4
B48.16=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O h5
B48.17=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O b5
B48.18=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Bd6
B48.19=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Ne5
B48.20=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Ne5 9.h3
B48.21=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Ne5 9.h3 Bc5
B48.22=Sicilianskt: Taimanov, 6.Be3 a6 7.Bd3 Nf6 8.O-O Ne5 9.h3 Bc5 10.Kh1
B49.1=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2
B49.2=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nge7
B49.3=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 b5
B49.4=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 b5 8.Nxc6
B49.5=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6
B49.6=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.a3
B49.7=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.a3 b5
B49.8=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.a3 Be7
B49.9=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.a3 Be7 9.O-O
B49.10=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O
B49.11=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O b5
B49.12=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Be7
B49.13=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4
B49.14=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Nxc6
B49.15=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4
B49.16=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4 O-O
B49.17=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4 Be7
B49.18=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4 Be7 10.Nxc6
B49.19=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4 Be7 10.Nxc6 bxc6
B49.20=Sicilianskt: Taimanov, 6.Be3 a6 7.Be2 Nf6 8.O-O Bb4 9.Na4 Be7 10.Nxc6 bxc6 11.Nb6
B50.1=Sicilianskt: 1.e4 c5 2.Nf3 d6
B50.2=Sicilianskt: Avb�jd vinggambit, 1.e4 c5 2.Nf3 d6 3.b4
B50.3=Sicilianskt: 2.Nf3 d6 3.b3
B50.4=Sicilianskt: 2.Nf3 d6 3.b3 e6
B50.5=Sicilianskt: 2.Nf3 d6 3.d3
B50.6=Sicilianskt: 2.Nf3 d6 3.g3
B50.7=Sicilianskt: 2.Nf3 d6 3.Bc4
B50.8=Sicilianskt: 2.Nf3 d6 3.Bc4 Nf6 4.d3
B50.9=Sicilianskt: 2.Nf3 d6 3.Nc3
B50.10=Sicilianskt: 2.Nf3 d6 3.Nc3 e6
B50.11=Sicilianskt: 2.Nf3 d6 3.Nc3 Nf6
B50.12=Sicilianskt: 2.Nf3 d6 3.c3
B50.13=Sicilianskt: 2.Nf3 d6 3.c3 Nf6
B50.14=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.h3
B50.15=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.h3 Nc6
B50.16=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Bc4
B50.17=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Bd3
B50.18=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Bd3 Nc6
B50.19=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Be2
B50.20=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Be2 Nc6
B50.21=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Be2 Nbd7
B50.22=Sicilianskt: 2.Nf3 d6 3.c3 Nf6 4.Be2 g6
B50.23=Sicilianskt: 2.Nf3 d6 3.c3, Torrevarianten
B51.1=Sicilianskt: 3.Bb5+
B51.2=Sicilianskt: 3.Bb5+ Nd7
B51.3=Sicilianskt: 3.Bb5+ Nd7 4.c3
B51.4=Sicilianskt: 3.Bb5+ Nd7 4.O-O
B51.5=Sicilianskt: 3.Bb5+ Nd7 4.O-O Nf6
B51.6=Sicilianskt: 3.Bb5+ Nd7 4.O-O Nf6 5.Re1 a6 6.Bf1
B51.7=Sicilianskt: 3.Bb5+ Nd7 4.d4
B51.8=Sicilianskt: 3.Bb5+ Nd7 4.d4 cxd4
B51.9=Sicilianskt: 3.Bb5+ Nd7 4.d4 Nf6
B51.10=Sicilianskt: 3.Bb5+ Nd7 4.d4 Nf6 5.Nc3
B51.11=Sicilianskt: 3.Bb5+ Nd7 4.d4 Nf6 5.Nc3 cxd4
B51.12=Sicilianskt: 3.Bb5+ Nd7 4.d4 Nf6 5.Nc3 cxd4 6.Qxd4
B51.13=Sicilianskt: 3.Bb5+ Nc6
B51.14=Sicilianskt: 3.Bb5+ Nc6 4.Bxc6+
B51.15=Sicilianskt: 3.Bb5+ Nc6 4.O-O
B51.16=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7
B51.17=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1
B51.18=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 a6
B51.19=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 Nf6
B51.20=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 Nf6 6.c3
B51.21=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 Nf6 6.c3 a6 7.Ba4
B51.22=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 Nf6 6.c3 a6 7.Bf1
B51.23=Sicilianskt: 3.Bb5+ Nc6 4.O-O Bd7 5.Re1 Nf6 6.c3 a6 7.Bf1 Bg4 8.h3
B52.1=Sicilianskt: 3.Bb5+ Bd7
B52.2=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Nxd7
B52.3=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Nxd7 5.O-O
B52.4=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Nxd7 5.O-O Ngf6
B52.5=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Nxd7 5.O-O Ngf6 6.Qe2
B52.6=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7
B52.7=Sicilianskt: 3.Bb5+, Sokolskyvarianten
B52.8=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6
B52.9=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6 6.O-O
B52.10=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6 6.O-O Nf6
B52.11=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6 6.Nc3
B52.12=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6 6.Nc3 Nf6
B52.13=Sicilianskt: 3.Bb5+, Sokolsky, 5...Nc6 6.Nc3 Nf6 7.O-O
B52.14=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O
B52.15=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6
B52.16=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6 6.Re1
B52.17=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6 6.Re1 Nf6
B52.18=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6 6.c3
B52.19=Sicilianskt: 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6 6.c3 Nf6
B52.20=Sicilianskt: Bronsteins gambit, 3.Bb5+ Bd7 4.Bxd7+ Qxd7 5.O-O Nc6 6.c3 Nf6 7.d4
B53.1=Sicilianskt: 1.e4 c5 2.Nf3 d6 3.d4
B53.2=Sicilianskt: 2...d6 3.d4 Nf6
B53.3=Sicilianskt: 2...d6 3.d4 cxd4
B53.4=Sicilianskt, Chekhovervarianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Qxd4
B53.5=Sicilianskt, Chekhover, 4...Bd7
B53.6=Sicilianskt, Chekhover, 4...a6
B53.7=Sicilianskt, Chekhover, 4...a6 5.Be3
B53.8=Sicilianskt, Chekhover, 4...a6 5.c4
B53.9=Sicilianskt, Chekhover, 4...a6 5.c4 Nc6 6.Qd2
B53.10=Sicilianskt, Chekhover, 4...a6 5.c4 Nc6 6.Qd2 g6
B53.11=Sicilianskt, Chekhover, 4...Nf6
B53.12=Sicilianskt, Chekhover, 4...Nf6 5.Nc3
B53.13=Sicilianskt, Chekhover, 4...Nc6
B53.14=Sicilianskt: Chekhover, Zaitsevvarianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Qxd4 Nc6 5.Bb5 Qd7
B53.15=Sicilianskt, Chekhover, 4...Nc6 5.Bb5 Bd7
B53.16=Sicilianskt, Chekhover, 4...Nc6 5.Bb5 Bd7 6.Bxc6 Bxc6
B53.17=Sicilianskt, Chekhover, 7.c4
B53.18=Sicilianskt, Chekhover, 7.c4 Nf6 8.Nc3 g6
B53.19=Sicilianskt, Chekhover, 7.Nc3
B53.20=Sicilianskt, Chekhover, 7.Nc3 Nf6 8.Bg5
B53.21=Sicilianskt, Chekhover, 7.Nc3 Nf6 8.Bg5 e6
B53.22=Sicilianskt, Chekhover, Huvudvarianten, 10.Qd3
B53.23=Sicilianskt, Chekhover, Huvudvarianten, 10.Rhe1
B53.24=Sicilianskt, Chekhover, Huvudvarianten, 10.Rhe1 O-O
B53.25=Sicilianskt, Chekhover, Huvudvarianten, 11.Qd2
B54.1=Sicilianskt: �ppet, 2...d6
B54.2=Sicilianskt: �ppet, 2...d6, 4...e5
B54.3=Sicilianskt: �ppet, 2...d6, 4...a6
B54.4=Sicilianskt: �ppet, 2...d6, 4...Nf6
B54.5=Sicilianskt: �ppet, 2...d6, 4...Nf6 5.Bd3
B54.6=Sicilianskt: Prins (Moskva)varianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.f3
B54.7=Sicilianskt: Prins (Moskva), 5...e6
B54.8=Sicilianskt: Prins (Moskva), 5...a6
B54.9=Sicilianskt: Prins (Moskva), 5...Nc6
B54.10=Sicilianskt: Prins (Moskva), 5...Nc6 6.c4 Nxd4
B54.11=Sicilianskt: Prins (Moskva), 5...Nc6 6.c4 Qb6
B54.12=Sicilianskt: Prins (Moskva), 5...e5
B54.13=Sicilianskt: Prins (Moskva), 5...e5 6.Nb3
B54.14=Sicilianskt: Prins (Moskva), 5...e5 6.Nb3 Be6
B54.15=Sicilianskt: Prins (Moskva), 5...e5 6.Nb3 d5
B55.1=Sicilianskt: Prins, Venice attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.f3 e5 6.Bb5+
B55.2=Sicilianskt: Prins, Venice attack, 6...Bd7
B55.3=Sicilianskt: Prins, Venice attack, 6...Nbd7
B55.4=Sicilianskt: Prins, Venice attack, 6...Nbd7 7.Nf5
B55.5=Sicilianskt: Prins, Venice attack, 6...Nbd7 7.Nf5 d5
B56.1=Sicilianskt: �ppet, 2...d6, 5.Nc3
B56.2=Sicilianskt: �ppet, 2...d6, 5.Nc3 e5
B56.3=Sicilianskt: Venice attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e5 6.Bb5+
B56.4=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nbd7
B56.5=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nbd7 6.Bc4
B56.6=Sicilianskt: �ppet, 2...d6, 5.Nc3 Bd7
B56.7=Sicilianskt: �ppet, 2...d6, 5.Nc3 Bd7 6.Bg5
B56.8=Sicilianskt: �ppet, 2...d6 5.Nc3 Nc6
B56.9=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.h3
B56.10=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.g3
B56.11=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.f4
B56.12=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.f3
B56.13=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.f3 e5
B56.14=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.f3 e5 7.Nb3
B56.15=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.f3 e5 7.Nb3 Be7
B56.16=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.Be3
B56.17=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.Be3 e5
B56.18=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.Be3 Ng4
B56.19=Sicilianskt: �ppet, 2...d6, 5.Nc3 Nc6 6.Be3 Ng4 7.Bb5
B57.1=Sicilianskt: Sozin, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Nc6 6.Bc4
B57.2=Sicilianskt: Sozin, Magnus Smiths f�lla, 6.Bc4 g6 7.Nxc6 bxc6 8.e5
B57.3=Sicilianskt: Sozin, 6...Bd7
B57.4=Sicilianskt: Sozin, 6...Bd7 7.O-O
B57.5=Sicilianskt: Sozin, Benkovarianten, 6.Bc4 Qb6
B57.6=Sicilianskt: Sozin, Benko, 7.Nde2
B57.7=Sicilianskt: Sozin, Benko, 7.Ndb5
B57.8=Sicilianskt: Sozin, Benko, 7.Nxc6
B57.9=Sicilianskt: Sozin, Benko, 7.Nxc6 bxc6 8.O-O g6
B57.10=Sicilianskt: Sozin, Benko, 7.Nb3
B57.11=Sicilianskt: Sozin, Benko, 7.Nb3 e6
B57.12=Sicilianskt: Sozin, Benko, 7.Nb3 e6 8.Be3
B57.13=Sicilianskt: Sozin, Benko, 7.Nb3 e6 8.Bf4
B57.14=Sicilianskt: Sozin, Benko, 7.Nb3 e6 8.O-O
B57.15=Sicilianskt: Sozin, Benko, 7.Nb3 e6 8.O-O Be7
B57.16=Sicilianskt: Sozin, Benko, 7.Nb3 e6 8.O-O Be7 9.Be3
B58.1=Sicilianskt: BoleSlaviskskyvarianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Nc6 6.Be2
B58.2=Sicilianskt: BoleSlavisksky, 6...Bd7
B58.3=Sicilianskt: BoleSlavisksky, 6...a6
B58.4=Sicilianskt: BoleSlavisksky, 6...Nxd4
B58.5=Sicilianskt: BoleSlavisksky, 6...e5
B58.6=Sicilianskt: BoleSlavisksky, 7.Ndb5
B58.7=Sicilianskt: BoleSlavisksky, Loumavarianten, 6.Be2 e5 7.Nxc6
B58.8=Sicilianskt: BoleSlavisksky, Loumavarianten, 6.Be2 e5 7.Nxc6 bxc6
B58.9=Sicilianskt: BoleSlavisksky, 7.Nf3
B58.10=Sicilianskt: BoleSlavisksky, 7.Nf3 h6
B58.11=Sicilianskt: BoleSlavisksky, 7.Nf3 h6 8.O-O
B58.12=Sicilianskt: BoleSlavisksky, 7.Nf3 h6 8.O-O Be7
B58.13=Sicilianskt: BoleSlavisksky, 7.Nf3 h6 8.O-O Be7 9.h3
B58.14=Sicilianskt: BoleSlavisksky, 7.Nf3 h6 8.O-O Be7 9.Re1
B58.15=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3
B58.16=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3 a6
B58.17=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3 Be6
B58.18=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3 Be6 11.Bf1
B58.19=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3 Be6 11.Bf1 Nb8
B58.20=Sicilianskt: BoleSlavisksky, 7.Nf3, 9.Re1 O-O 10.h3 Be6 11.Bf1 Nb8 12.b3
B59.1=Sicilianskt: BoleSlavisksky, 7.Nb3
B59.2=Sicilianskt: BoleSlavisksky, 7.Nb3 Be6
B59.3=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7
B59.4=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.Bg5
B59.5=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.Be3
B59.6=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O
B59.7=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O
B59.8=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.Bg5
B59.9=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.Kh1
B59.10=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.f4
B59.11=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.Be3
B59.12=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.Be3 Be6
B59.13=Sicilianskt: BoleSlavisksky, 7.Nb3 Be7 8.O-O O-O 9.Be3 a5
B60.1=Sicilianskt: Richter-Rauzer, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Nc6 6.Bg5
B60.2=Sicilianskt: Richter-Rauzer, Bondarevskyvarianten, 6.Bg5 g6
B60.3=Sicilianskt: Richter-Rauzer, 6...Qa5
B60.4=Sicilianskt: Richter-Rauzer, 6...Qb6
B60.5=Sicilianskt: Richter-Rauzer, 6...a6
B60.6=Sicilianskt: Richter-Rauzer, Larsenvarianten, 6.Bg5 Bd7
B60.7=Sicilianskt: Richter-Rauzer, Larsen, 7.Nb3
B60.8=Sicilianskt: Richter-Rauzer, Larsen, 7.Bxf6
B60.9=Sicilianskt: Richter-Rauzer, Larsen, 7.Be2
B60.10=Sicilianskt: Richter-Rauzer, Larsen, 7.Be2 a6
B60.11=Sicilianskt: Richter-Rauzer, Larsen, 7.Be2 Qa5
B61.1=Sicilianskt: Richter-Rauzer, Larsen, 7.Qd2
B61.2=Sicilianskt: Richter-Rauzer, Larsen, 7.Qd2 a6
B61.3=Sicilianskt: Richter-Rauzer, Larsen, 7.Qd2 Nxd4
B61.4=Sicilianskt: Richter-Rauzer, Larsen, 7.Qd2 Rc8
B61.5=Sicilianskt: Richter-Rauzer, Larsen, 7.Qd2 Rc8 8.O-O-O
B62.1=Sicilianskt: Richter-Rauzer, 6...e6
B62.2=Sicilianskt: Richter-Rauzer, 6...e6 7.Be2
B62.3=Sicilianskt: Richter-Rauzer, Podebradyvarianten, 6...e6 7.Nb3
B62.4=Sicilianskt: Richter-Rauzer, Richter attack, 6...e6 7.Nxc6
B62.5=Sicilianskt: Richter-Rauzer, Keresvarianten, 6...e6 7.Qd3
B62.6=Sicilianskt: Richter-Rauzer, Margate (Alekhine)varianten, 6...e6 7.Bb5
B62.7=Sicilianskt: Richter-Rauzer, Margate (Alekhine)varianten, 7...Bd7
B63.1=Sicilianskt: Richter-Rauzer, Rauzer attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 Nc6 6.Bg5 e6 7.Qd2
B63.2=Sicilianskt: Richter-Rauzer, 7.Qd2 Nxd4
B63.3=Sicilianskt: Richter-Rauzer, 7.Qd2 Qb6
B63.4=Sicilianskt: Richter-Rauzer, 7.Qd2 Qb6 8.Nb3
B63.5=Sicilianskt: Richter-Rauzer, 7.Qd2 Qb6 8.Nb3 a6
B63.6=Sicilianskt: Richter-Rauzer, 7.Qd2 Qb6 8.Nb3 a6 9.O-O-O
B63.7=Sicilianskt: Richter-Rauzer, 7.Qd2 Qb6 8.Nb3 a6 9.O-O-O Be7
B63.8=Sicilianskt: Richter-Rauzer, 7.Qd2 h6
B63.9=Sicilianskt: Richter-Rauzer, 7.Qd2 h6 8.Bxf6 gxf6 9.O-O-O a6
B63.10=Sicilianskt: Richter-Rauzer, 7.Qd2 h6 8.Bxf6 gxf6 9.O-O-O a6 10.f4
B63.11=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7
B63.12=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O
B63.13=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O Nxd4
B63.14=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O Nxd4
B63.15=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O Nxd4 9.Qxd4 O-O
B63.16=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O
B63.17=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7, 9.f3
B63.18=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7, 9.Nb3
B63.19=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7, 9.Nb3 a5
B63.20=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7, 9.Nb3 a6
B63.21=Sicilianskt: Richter-Rauzer, Podebradvarianten, 7.Qd2 Be7 8.O-O-O O-O 9.Nb3 Qb6
B63.22=Sicilianskt: Richter-Rauzer, Podebradvarianten, 10.f3
B63.23=Sicilianskt: Richter-Rauzer, Podebradvarianten, 10.f3 Rd8
B63.24=Sicilianskt: Richter-Rauzer, Podebradvarianten, 10.f3 Rd8 11.Kb1
B64.1=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4
B64.2=Sicilianskt: Richter-Rauzer, Gellervarianten, 7.Qd2 Be7 8.O-O-O O-O 9.f4 e5
B64.3=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7, 9.f4 h6
B64.4=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 h6 10.Bh4 Bd7
B65.1=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4
B65.2=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4 10.Qxd4
B65.3=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4 10.Qxd4 h6
B65.4=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4 10.Qxd4 Qa5
B65.5=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4 10.Qxd4 Qa5 11.Kb1
B65.6=Sicilianskt: Richter-Rauzer, 7.Qd2 Be7 8.O-O-O O-O 9.f4 Nxd4 10.Qxd4 Qa5 11.Bc4
B66.1=Sicilianskt: Richter-Rauzer, 7...a6
B66.2=Sicilianskt: Richter-Rauzer, 7...a6 8.Be2
B66.3=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O
B66.4=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O Be7
B66.5=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O Nxd4
B66.6=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O Nxd4 9.Qxd4
B66.7=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O Nxd4 9.Qxd4 Be7
B66.8=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6
B66.9=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Bf4
B66.10=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Bf4, 11.f3
B66.11=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3
B66.12=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Qc7
B66.13=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Bd7
B66.14=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Bd7 10.f3
B66.15=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7
B66.16=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7 10.f3
B66.17=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7 10.f3 Nxd4
B66.18=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7 10.f3 Nxd4 11.Bxd4
B66.19=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7 10.f4
B66.20=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O h6 9.Be3 Be7 10.f4 Nxd4
B67.1=Sicilianskt: Richter-Rauzer, 7...a6 8.O-O-O Bd7
B67.2=Sicilianskt: Richter-Rauzer, 7...a6, 9.Be2
B67.3=Sicilianskt: Richter-Rauzer, 7...a6, 9.f3
B67.4=Sicilianskt: Richter-Rauzer, 7...a6, 9.f3 Rc8
B67.5=Sicilianskt: Richter-Rauzer, 7...a6, 9.f3 Be7
B67.6=Sicilianskt: Richter-Rauzer, 7...a6, 9.f3 Be7 10.h4
B67.7=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4
B67.8=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 h6
B67.9=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 h6 10.Bh4
B67.10=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 h6 10.Bh4 g5
B67.11=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5
B67.12=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Nxc6
B67.13=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6
B67.14=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6
B67.15=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.f5
B67.16=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.Nxc6
B67.17=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.Nxc6 Bxc6 12.Qe1
B67.18=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.Kb1
B67.19=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.Kb1 Qb6
B67.20=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 b5 10.Bxf6 gxf6 11.Kb1 Qb6 12.Nxc6
B68.1=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7
B68.2=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Be2
B68.3=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Be2 Qc7
B68.4=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3
B68.5=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5
B68.6=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5 11.e5
B69.1=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5 11.Bxf6
B69.2=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5 11.Bxf6 gxf6
B69.3=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5 11.Bxf6 gxf6 12.Kb1
B69.4=Sicilianskt: Richter-Rauzer, 7...a6, 9.f4 Be7 10.Nf3 b5 11.Bxf6 gxf6 12.f5
B70.1=Sicilianskt: Draken, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 g6
B70.2=Sicilianskt: Draken, 6.f3
B70.3=Sicilianskt: Draken, 6.g3
B70.4=Sicilianskt: Draken, 6.g3 Nc6
B70.5=Sicilianskt: Draken, 6.g3 Nc6 7.Bg2
B70.6=Sicilianskt: Draken, 6.g3 Nc6 7.Nde2
B70.7=Sicilianskt: Draken, 6.Bg5
B70.8=Sicilianskt: Draken, 6.Bg5
B70.9=Sicilianskt: Draken, 6.Bc4
B70.10=Sicilianskt: Draken, 6.Bc4 Bg7
B70.11=Sicilianskt: Draken, 6.Bc4 Bg7 7.h3
B70.12=Sicilianskt: Draken, 6.Bc4 Bg7 7.O-O
B70.13=Sicilianskt: Draken, 6.Be2
B70.14=Sicilianskt: Draken, 6.Be2 Nc6
B70.15=Sicilianskt: Draken, 6.Be2 a6
B70.16=Sicilianskt: Draken, 6.Be2 a6 7.a4 Bg7
B70.17=Sicilianskt: Draken, 6.Be2 Bg7
B70.18=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O
B70.19=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O Nc6
B70.20=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O Nc6 8.Nb3
B70.21=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O Nc6 8.Nb3 O-O
B70.22=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O
B70.23=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Re1
B70.24=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Re1 Nc6
B70.25=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Re1 Nc6 9.Nb3
B70.26=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Re1 Nc6 9.Nb3 Be6
B70.27=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5
B70.28=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5
B70.29=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5 Nc6 9.Nb3
B70.30=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5 Nc6 9.Nb3 a6
B70.31=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5 Nc6 9.Nb3 Be6
B70.32=Sicilianskt: Draken, 6.Be2 Bg7 7.O-O O-O 8.Bg5 Nc6 9.Nb3 Be6 10.Kh1
B71.1=Sicilianskt: Draken, Levenfishvarianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 g6 6.f4
B71.2=Sicilianskt: Draken, Levenfish, 6...Bg7
B71.3=Sicilianskt: Draken, Levenfish, 6...Bg7 7.e5
B71.4=Sicilianskt: Draken, Levenfish, 6...Nbd7
B71.5=Sicilianskt: Draken, Levenfish, 6...Nc6
B71.6=Sicilianskt: Draken, Levenfish, 6...Nc6 7.Bb5
B71.7=Sicilianskt: Draken, Levenfish, 6...Nc6 7.Nf3
B71.8=Sicilianskt: Draken, Levenfish, 6...Nc6 7.Nxc6
B72.1=Sicilianskt: Draken, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 g6 6.Be3
B72.2=Sicilianskt: Draken, 6.Be3 Bg7
B72.3=Sicilianskt: Draken, 6.Be3 Bg7 7.Qd2
B72.4=Sicilianskt: Draken, 6.Be3 Bg7 7.Bc4
B72.5=Sicilianskt: Draken, 6.Be3 Bg7 7.Bc4 Nc6
B72.6=Sicilianskt: Draken, 6.Be3 Bg7 7.Bc4 O-O
B72.7=Sicilianskt: Draken, Klassisk attack, 6.Be3 Bg7 7.Be2
B72.8=Sicilianskt: Draken, Klassisk attack, 6.Be3 Bg7 7.Be2 O-O
B72.9=Sicilianskt: Draken, Klassisk attack, 6.Be3 Bg7 7.Be2 O-O 8.O-O
B72.10=Sicilianskt: Draken, Klassisk, Amsterdamvarianten, 6.Be3 Bg7 7.Be2 Nc6 8.Qd2
B72.11=Sicilianskt: Draken, Klassisk, Grigorievvarianten, 6.Be3 Bg7 7.Be2 Nc6 8.Qd2 O-O 9.O-O-O
B72.12=Sicilianskt: Draken, Klassisk, Nottinghamvarianten, 6.Be3 Bg7 7.Be2 Nc6 8.Nb3
B73.1=Sicilianskt: Draken, Klassisk, 8.O-O
B73.2=Sicilianskt: Draken, Klassisk, 8.O-O O-O
B73.3=Sicilianskt: Draken, Klassisk, 9.Kh1
B73.4=Sicilianskt: Draken, Klassisk, Richtervarianten, 8.O-O O-O 9.Qd2
B73.5=Sicilianskt: Draken, Klassisk, 9.f4
B73.6=Sicilianskt: Draken, Klassisk, Zollner gambit, 8.O-O O-O 9.f4 Qb6 10.e5
B74.1=Sicilianskt: Draken, Klassisk, 9.Nb3
B74.2=Sicilianskt: Draken, Klassisk, 9.Nb3 b6
B74.3=Sicilianskt: Draken, Klassisk, Alekhinevarianten, 9.Nb3 a5
B74.4=Sicilianskt: Draken, Klassisk, 9.Nb3 a6
B74.5=Sicilianskt: Draken, Klassisk, 9.Nb3 Be6
B74.6=Sicilianskt: Draken, Klassisk, 9.Nb3 Be6 10.f4
B74.7=Sicilianskt: Draken, Klassisk, 9.Nb3 Be6 10.f4 Rc8
B74.8=Sicilianskt: Draken, Klassisk, Tartakowervarianten, 9.Nb3 Be6 10.f4 Qc8
B74.9=Sicilianskt: Draken, Klassisk, Maroczyvarianten, 9.Nb3 Be6 10.f4 Na5
B74.10=Sicilianskt: Draken, Klassisk, Stockholmattacken, 9.Nb3 Be6 10.f4 Na5 11.f5 Bc4 12.Nxa5 Bxe2 13.Qxe2 Qxa5 14.g4
B74.11=Sicilianskt: Draken, Klassisk, Spielmannvarianten, 9.Nb3 Be6 10.f4 Na5 11.f5 Bc4 12.Bd3
B74.12=Sicilianskt: Draken, Klassisk, Bernards f�rsvar, 9.Nb3 Be6 10.f4 Na5 11.f5 Bc4 12.Bd3 Bxd3 13.cxd3 d5
B75.1=Sicilianskt: Draken, Jugoslavisk attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 g6 6.Be3 Bg7 7.f3
B75.2=Sicilianskt: Draken, Jugoslavisk, 7...a6
B75.3=Sicilianskt: Draken, Jugoslavisk, 7...Nc6
B75.4=Sicilianskt: Draken, Jugoslavisk, 7...Nc6 8.Bc4
B75.5=Sicilianskt: Draken, Jugoslavisk, 7...Nc6 8.Qd2
B75.6=Sicilianskt: Draken, Jugoslavisk, 7...Nc6 8.Qd2 Bd7
B75.7=Sicilianskt: Draken, Jugoslavisk, 7...Nc6 8.Qd2 Bd7 9.O-O-O
B75.8=Sicilianskt: Draken, Jugoslavisk, 7...Nc6 8.Qd2 Bd7 9.O-O-O Rc8
B76.1=Sicilianskt: Draken, Jugoslavisk, 7.f3 O-O
B76.2=Sicilianskt: Draken, Jugoslavisk, 7.f3 O-O 8.Qd2
B76.3=Sicilianskt: Draken, Jugoslavisk, 8.Qd2 Nc6
B76.4=Sicilianskt: Draken, Jugoslavisk, 9.g4
B76.5=Sicilianskt: Draken, Jugoslavisk, 9.g4 Be6
B76.6=Sicilianskt: Draken, Jugoslavisk, 9.g4 Nxd4
B76.7=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O
B76.8=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Bd7
B76.9=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Bd7 10.g4
B76.10=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Nxd4
B76.11=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Nxd4 10.Bxd4 Be6
B76.12=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Nxd4: 11.Kb1
B76.13=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Nxd4: 11.Kb1 Qc7
B76.14=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O Nxd4: 11.Kb1 Qc7 12.g4
B76.15=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5
B76.16=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5 10.Qe1
B76.17=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5 10.exd5
B76.18=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5 10.exd5 Nxd5 11.Nxc6
B76.19=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5: 12.Nxd5
B76.20=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5: 12.Bd4
B76.21=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5: 12.Bd4 e5
B76.22=Sicilianskt: Draken, Jugoslavisk, 9.O-O-O d5: 12.Bd4 e5 13.Bc5 Be6
B77.1=Sicilianskt: Draken, Jugoslavisk, 9.Bc4
B77.2=Sicilianskt: Draken, Jugoslavisk, Byrnevarianten, 9.Bc4 a5
B77.3=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Ne5
B77.4=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Nd7
B77.5=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Nxd4
B77.6=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Bd7
B77.7=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Bd7 10.Bb3
B77.8=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Bd7 10.g4
B77.9=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Bd7 10.h4
B77.10=Sicilianskt: Draken, Jugoslavisk, 9.Bc4 Bd7 10.h4 Rc8
B78.1=Sicilianskt: Draken, Jugoslavisk, 10.O-O-O
B78.2=Sicilianskt: Draken, Jugoslavisk, 10.O-O-O Ne5
B78.3=Sicilianskt: Draken, Jugoslavisk, 10.O-O-O Rc8
B78.4=Sicilianskt: Draken, Jugoslavisk, 10.O-O-O Rc8 11.Bb3
B78.5=Sicilianskt: Draken, Jugoslavisk, Moderna Huvudvarianten, 10.O-O-O Rc8 11.Bb3 Ne5
B78.6=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.Kb1
B78.7=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.Kb1
B78.8=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.Kb1: 14.g4 b5
B78.9=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4
B78.10=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 Nc4
B78.11=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 Nc4: 14.g4
B78.12=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 Nc4: 14.h5
B78.13=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5
B78.14=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Kb1
B78.15=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bh6
B78.16=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bh6 Bxh6
B78.17=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bg5
B78.18=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bg5 Rc5
B78.19=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bg5 Rc5 14.g4
B78.20=Sicilianskt: Draken, Jugoslavisk, Huvudvarianten, 12.h4 h5 13.Bg5 Rc5 14.Kb1
B78.21=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 10.O-O-O Qa5
B78.22=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 11.Bb3 Rac8
B78.23=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 11.Bb3 Rfc8
B79.1=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4
B79.2=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 h5
B79.3=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 Ne5
B79.4=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 Ne5 13.Kb1
B79.5=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 Ne5 13.Kb1 Nc4
B79.6=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 Ne5 13.g4
B79.7=Sicilianskt: Draken, Jugoslavisk, Gamla Huvudvarianten, 12.h4 Ne5 13.h5
B80.1=Sicilianskt: Scheveningen, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6
B80.2=Sicilianskt: Scheveningen, 6.Be3
B80.3=Sicilianskt: Scheveningen, 6.Be3 Nc6
B80.4=Sicilianskt: Scheveningen, 6.Be3 Nc6
B80.5=Sicilianskt: Scheveningen, 6.Be3 a6
B80.6=Sicilianskt: Scheveningen, 7.Qd2
B80.7=Sicilianskt: Scheveningen, Engelsk attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Be3 a6 7.f3
B80.8=Sicilianskt: Scheveningen, Engelsk attack, 7...Nc6
B80.9=Sicilianskt: Scheveningen, Engelsk, 7...Nc6 8.Qd2
B80.10=Sicilianskt: Scheveningen, Engelsk, 7...Nc6 8.Qd2
B80.11=Sicilianskt: Scheveningen, Engelsk attack, 7...b5
B80.12=Sicilianskt: Scheveningen, Engelsk, 7...b5 8.Qd2
B80.13=Sicilianskt: Scheveningen, Engelsk, 7...b5, 8.Qd2 Bb7
B80.14=Sicilianskt: Scheveningen, Engelsk, 7...b5 8.Qd2 Bb7
B80.15=Sicilianskt: Scheveningen, Engelsk, 7...b5 8.Qd2 Nbd7
B80.16=Sicilianskt: Scheveningen, Vitolinvarianten, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Bb5+
B80.17=Sicilianskt: Scheveningen, Vitolins, 6...Bd7
B80.18=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3
B80.19=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 a6
B80.20=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6
B80.21=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 a6
B80.22=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 a6 8.O-O
B80.23=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 a6 8.O-O Bd7
B80.24=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 Qc7
B80.25=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 Qc7 8.O-O a6
B80.26=Sicilianskt: Scheveningen, Fianchettovarianten, 6.g3 Nc6 7.Bg2 Qc7 8.O-O a6 9.Re1 Be7
B81.1=Sicilianskt: Scheveningen, Keres attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.g4
B81.2=Sicilianskt: Scheveningen, Keres, 6...e5
B81.3=Sicilianskt: Scheveningen, Keres, 6...a6
B81.4=Sicilianskt: Scheveningen, Keres, Perenyi attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.g4 a6 7.Be3
B81.5=Sicilianskt: Scheveningen, Keres, Perenyi attack, 7...e5
B81.6=Sicilianskt: Scheveningen, Keres, Perenyi attack, 7...h6
B81.7=Sicilianskt: Scheveningen, Keres, Perenyi attack, 7...h6 8.f4
B81.8=Sicilianskt: Scheveningen, Keres, 6...h6
B81.9=Sicilianskt: Scheveningen, Keres, 6...h6 7.h3 Nc6 8.Bg2
B81.10=Sicilianskt: Scheveningen, Keres, 6...h6 7.h3 Nc6 8.Bg2
B81.11=Sicilianskt: Scheveningen, Keres, 6...h6 7.h3 a6 8.Bg2
B81.12=Sicilianskt: Scheveningen, Keres, 6...h6 7.h4
B81.13=Sicilianskt: Scheveningen, Keres, 6...h6 7.h4 Be7
B81.14=Sicilianskt: Scheveningen, Keres, 6...h6 7.h4 Nc6
B81.15=Sicilianskt: Scheveningen, Keres, 6...h6 7.h4 Nc6 8.Rg1
B81.16=Sicilianskt: Scheveningen, Keres, 6...h6 7.h4 Nc6 8.Rg1 h5
B81.17=Sicilianskt: Scheveningen, Keres, 6...h6 7.g5
B81.18=Sicilianskt: Scheveningen, Keres, 6...h6 7.Rg1
B81.19=Sicilianskt: Scheveningen, Keres, 6...Nc6
B81.20=Sicilianskt: Scheveningen, Keres, 6...Nc6 7.g5 Nd7
B81.21=Sicilianskt: Scheveningen, Keres, 6...Nc6 7.g5 Nd7 8.Be3
B81.22=Sicilianskt: Scheveningen, Keres, 6...Nc6 7.g5 Nd7 8.Be3 Be7
B82.1=Sicilianskt: Scheveningen, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.f4
B82.2=Sicilianskt: Scheveningen, 6.f4 Qb6
B82.3=Sicilianskt: Scheveningen, 6.f4 Be7
B82.4=Sicilianskt: Scheveningen, 6.f4 a6
B82.5=Sicilianskt: Scheveningen, 6.f4 a6 7.Be3
B82.6=Sicilianskt: Scheveningen, 6.f4 a6 7.Be3 b5
B82.7=Sicilianskt: Scheveningen, 6.f4 Nc6
B82.8=Sicilianskt: Scheveningen, 6.f4 Nc6 7.Be3
B82.9=Sicilianskt: Scheveningen, 6.f4 Nc6 7.Be3 Qc7
B82.10=Sicilianskt: Scheveningen, 6.f4 Nc6 7.Be3 Be7
B82.11=Sicilianskt: Scheveningen, Talvarianten, 6.f4 Nc6 7.Be3 Be7 8.Qf3
B82.12=Sicilianskt: Scheveningen, Talvarianten, 8...e5
B82.13=Sicilianskt: Scheveningen, Talvarianten, 8...Qc7
B83.1=Sicilianskt: Scheveningen, 6.Be2
B83.2=Sicilianskt: Scheveningen, 6.Be2
B83.3=Sicilianskt: Scheveningen, Moderna, 6.Be2 Nc6
B83.4=Sicilianskt: Scheveningen, Moderna, 6.Be2 Nc6 7.O-O Be7
B83.5=Sicilianskt: Scheveningen, Moderna, 6.Be2 Nc6 7.O-O Be7 8.Be3 O-O
B83.6=Sicilianskt: Scheveningen, Moderna, 9.f4
B83.7=Sicilianskt: Scheveningen, Moderna, 9.f4 e5
B83.8=Sicilianskt: Scheveningen, Moderna, 9.f4 e5 10.Nb3
B83.9=Sicilianskt: Scheveningen, Moderna, 9.f4 e5 10.Nb3 exf4 11.Bxf4
B83.10=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7
B83.11=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7 10.Nb3
B83.12=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7 10.Nb3 a6
B83.13=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7 10.Nb3 a6 11.a4
B83.14=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7 10.Kh1
B83.15=Sicilianskt: Scheveningen, Moderna, 9.f4 Bd7 10.Qe1
B84.1=Sicilianskt: Scheveningen, Klassisk, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Be2 a6
B84.2=Sicilianskt: Scheveningen, Klassisk, 7.a4
B84.3=Sicilianskt: Scheveningen, Klassisk, 7.f4
B84.4=Sicilianskt: Scheveningen, Klassisk, 7.Be3
B84.5=Sicilianskt: Scheveningen, Klassisk, 7.O-O
B84.6=Sicilianskt: Scheveningen, Klassisk, 7.O-O Nbd7
B84.7=Sicilianskt: Scheveningen, Klassisk, 7.O-O Nbd7 8.a4
B84.8=Sicilianskt: Scheveningen, Klassisk, 7.O-O Nbd7 8.f4
B84.10=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7
B84.11=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.Kh1
B84.12=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.Kh1 Nc6
B84.13=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.a4
B84.14=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.a4 Nc6
B84.15=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.Bf3
B84.16=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.Be3
B84.17=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.Be3 Nc6
B84.18=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.f4
B84.19=Sicilianskt: Scheveningen, Klassisk, 7.O-O Qc7 8.f4 Nc6
B84.20=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7
B84.21=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7 8.f4
B84.22=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7 8.f4 Qc7
B84.23=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7 8.f4 Qc7 9.Be3
B84.25=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7 8.f4 Qc7 9.Kh1
B85.1=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9.Be3
B85.3=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6
B85.4=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Qe1
B85.5=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Qe1 Qc7
B85.6=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Qe1 Qc7 11.Qg3
B85.7=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Kh1
B85.8=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Kh1 Bd7
B85.9=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.Kh1 Qc7
B85.10=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.a4
B85.11=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.a4 Bd7
B85.12=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.a4 Qc7
B85.13=Sicilianskt: Scheveningen, Klassisk, Huvudvarianten, 9...Nc6 10.a4 Qc7 11.Kh1
B84.26=Sicilianskt: Scheveningen, Klassisk, 7.O-O Be7 8.f4 O-O
B86.1=Sicilianskt: Sozin-Scheveningen, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Bc4
B86.2=Sicilianskt: Sozin-Scheveningen, 6...Qb6
B86.3=Sicilianskt: Sozin-Najdorf
B86.4=Sicilianskt: Sozin-Najdorf, 7.Bb3
B86.5=Sicilianskt: Sozin-Najdorf, 7.Bb3 Be7
B87.1=Sicilianskt: Sozin-Najdorf, 7.Bb3 b5
B87.2=Sicilianskt: Sozin-Najdorf, 7.Bb3 b5 8.O-O
B87.3=Sicilianskt: Sozin-Najdorf, 7.Bb3 b5 8.O-O Be7
B87.4=Sicilianskt: Sozin-Najdorf, 7.Bb3 b5 8.O-O Be7 9.Qf3
B87.5=Sicilianskt: Sozin-Najdorf, 7.Bb3 b5 8.O-O Be7 9.f4
B88.1=Sicilianskt: Sozin-Scheveningen, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Bc4 Nc6
B88.2=Sicilianskt: Sozin-Scheveningen, 7.O-O
B88.3=Sicilianskt: Sozin-Scheveningen, 7.Bb3
B88.4=Sicilianskt: Sozin-Scheveningen, 7.Bb3
B88.5=Sicilianskt: Sozin, Fischervarianten, 6.Bc4 Nc6 7.Bb3 Be7 8.Be3 O-O 9.f4
B89.1=Sicilianskt: Sozin, 7.Be3
B89.2=Sicilianskt: Sozin, 7.Be3 a6
B89.3=Sicilianskt: Velimirovic mot 7...a6
B89.4=Sicilianskt: Sozin, 7.Be3 Be7
B89.5=Sicilianskt: Velimirovic, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 e6 6.Bc4 Nc6 7.Be3 Be7 8.Qe2
B89.6=Sicilianskt: Velimirovic, 9.O-O-O
B89.7=Sicilianskt: Velimirovic, 9.O-O-O Qc7
B89.8=Sicilianskt: Velimirovic, 9.O-O-O Qc7 10.Bb3 a6
B90.1=Sicilianskt: Najdorf, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 a6
B90.2=Sicilianskt: Najdorf, 6.a4
B90.3=Sicilianskt: Najdorf, 6.a4 e5
B90.4=Sicilianskt: Najdorf, 6.f3
B90.5=Sicilianskt: Najdorf, Adams attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 a6 6.h3
B90.6=Sicilianskt: Najdorf, Fischer-Sozin attack, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 a6 6.Bc4
B90.7=Sicilianskt: Najdorf, 6.Be3
B90.8=Sicilianskt: Najdorf, 6.Be3 Ng4
B90.9=Sicilianskt: Najdorf, 6.Be3 Ng4 7.Bg5
B90.10=Sicilianskt: Najdorf, 6.Be3 Ng4 7.Bg5 h6 8.Bh4 g5 9.Bg3 Bg7
B90.11=Sicilianskt: Najdorf, 6.Be3 Ng4 7.Bg5 h6 8.Bh4 g5 9.Bg3 Bg7 10.Be2
B90.12=Sicilianskt: Najdorf, 6.Be3 Ng4 7.Bg5 h6 8.Bh4 g5 9.Bg3 Bg7 10.Be2 h5
B90.13=Sicilianskt: Najdorf, 6.Be3 e5
B90.14=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3
B90.15=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.Qd2
B90.16=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3
B90.17=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7
B90.18=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7 9.Qd2
B90.19=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7 9.Qd2 Nbd7
B90.20=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7 9.Qd2 O-O
B90.21=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Nbd7
B90.22=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7 9.Qd2
B90.23=Sicilianskt: Najdorf, 6.Be3 e5 7.Nb3 Be6 8.f3 Be7 9.Qd2 b5
B91.1=Sicilianskt: Najdorf, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 a6 6.g3
B91.2=Sicilianskt: Najdorf, 6.g3 b5
B91.3=Sicilianskt: Najdorf, 6.g3 g6
B91.4=Sicilianskt: Najdorf, 6.g3 Nc6
B91.5=Sicilianskt: Najdorf, 6.g3 Bg4
B91.6=Sicilianskt: Najdorf, 6.g3 e5
B91.7=Sicilianskt: Najdorf, 6.g3 e5 7.Nb3
B91.8=Sicilianskt: Najdorf, 6.g3 e5 7.Nb3 Be7
B91.9=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2
B91.10=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2 b5
B91.11=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2 Nbd7
B91.12=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2 Be7
B91.13=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2 Be7 8.Bg2 Nbd7
B91.14=Sicilianskt: Najdorf, 6.g3 e5 7.Nde2 Be7 8.Bg2 O-O
B92.1=Sicilianskt: Najdorf, 6.Be2
B92.2=Sicilianskt: Najdorf, 6.Be2 Nbd7
B92.3=Sicilianskt: Najdorf, 6.Be2 e5
B92.4=Sicilianskt: Najdorf, 6.Be2 e5 7.Nf3
B92.5=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3
B92.6=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7
B92.7=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.Be3
B92.8=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.Be3 Be6
B92.9=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O
B92.10=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O Be6
B92.11=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O Be6 9.f4
B92.12=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O
B92.13=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Be3
B92.14=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Be3 Be6
B92.15=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Be3 Be6 10.a4
B92.16=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Be3 Be6 10.Nd5
B92.17=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Be3 Be6 10.Qd2
B92.18=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Kh1
B92.19=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Kh1 Be6
B92.20=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Kh1 Nc6
B92.21=Sicilianskt: Najdorf, 6.Be2 e5 7.Nb3 Be7 8.O-O O-O 9.Kh1 Qc7
B93.1=Sicilianskt: Najdorf, 6.f4
B93.2=Sicilianskt: Najdorf, 6.f4 Nc6
B93.3=Sicilianskt: Najdorf, 6.f4 Nbd7
B93.5=Sicilianskt: Najdorf, 6.f4 Qc7
B93.6=Sicilianskt: Najdorf, 6.f4 Qc7 7.Bd3
B93.7=Sicilianskt: Najdorf, 6.f4 Qc7 7.Bd3 g6
B93.8=Sicilianskt: Najdorf, 6.f4 Qc7 7.Nf3
B93.9=Sicilianskt: Najdorf, 6.f4 Qc7 7.Nf3 Nbd7
B93.10=Sicilianskt: Najdorf, 6.f4 Qc7 7.Nf3 Nbd7 8.Bd3
B93.11=Sicilianskt: Najdorf, 6.f4 e5
B93.12=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3
B93.13=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Qc7
B93.14=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Qc7 8.a4
B93.15=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7
B93.16=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.Bd3
B93.17=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4
B93.18=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Qc7
B93.19=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Be7
B93.20=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Be7 9.Bc4
B93.21=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Be7 9.Bd3
B93.22=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Be7 9.Bd3 O-O 10.O-O Nc5
B93.23=Sicilianskt: Najdorf, 6.f4 e5 7.Nf3 Nbd7 8.a4 Be7 9.Bd3 O-O 10.O-O exf4
B94.1=Sicilianskt: Najdorf, 6.Bg5
B94.2=Sicilianskt: Najdorf, 6.Bg5 b5
B94.3=Sicilianskt: Najdorf, 6.Bg5 e5
B94.4=Sicilianskt: Najdorf, 6.Bg5 Nbd7
B94.5=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.f4
B94.6=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.Bc4
B94.7=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.Bc4 e6
B94.8=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.Bc4 e6 8.O-O
B94.9=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.Bc4 Qa5
B94.10=Sicilianskt: Najdorf, 6.Bg5 Nbd7 7.Bc4 Qa5 8.Qd2 e6 9.O-O-O
B95.1=Sicilianskt: Najdorf, 6...e6
B95.2=Sicilianskt: Najdorf, 6...e6 7.Bd3
B95.3=Sicilianskt: Najdorf, 6...e6 7.Be2
B95.4=Sicilianskt: Najdorf, 6...e6 7.Qe2
B95.5=Sicilianskt: Najdorf, 6...e6 7.Qd2
B95.6=Sicilianskt: Najdorf, 6...e6 7.Qd2 Be7
B95.7=Sicilianskt: Najdorf, 6...e6 7.Qd2 Be7 8.O-O-O
B95.8=Sicilianskt: Najdorf, 6...e6 7.Qd3
B95.9=Sicilianskt: Najdorf, 6...e6 7.Qd3 Nc6
B95.10=Sicilianskt: Najdorf, 6...e6 7.Qf3
B95.11=Sicilianskt: Najdorf, 6...e6 7.Qf3 Nbd7
B95.12=Sicilianskt: Najdorf, 6...e6 7.Qf3 Be7
B95.13=Sicilianskt: Najdorf, 6...e6 7.Qf3 Be7 8.O-O-O Nbd7
B95.14=Sicilianskt: Najdorf, 6...e6 7.Qf3 h6
B96.1=Sicilianskt: Najdorf, 7.f4
B96.2=Sicilianskt: Najdorf, 7.f4 h6
B96.3=Sicilianskt: Najdorf, F�rdr�jd f�rgiftad bonde, 7.f4 h6 8.Bh4 Qb6
B96.4=Sicilianskt: Najdorf, 7.f4 Nc6
B96.5=Sicilianskt: Najdorf, 7.f4 Nc6 8.e5
B96.6=Sicilianskt: Najdorf, 7.f4 Nc6 8.Nxc6
B96.7=Sicilianskt: Najdorf, 7.f4 Bd7
B96.8=Sicilianskt: Najdorf, 7.f4 Qc7
B96.9=Sicilianskt: Najdorf, 7.f4 Qc7 8.Bxf6
B96.10=Sicilianskt: Najdorf, 7.f4 Qc7 8.Qf3
B96.11=Sicilianskt: Najdorf, 7.f4 Qc7 8.Qf3 b5
B96.12=Sicilianskt: Najdorf, 7.f4 Qc7 8.Qf3 b5 9.f5
B96.13=Sicilianskt: Najdorf, 7.f4 Qc7 8.Qf3 b5 9.O-O-O
B96.14=Sicilianskt: Najdorf, 7.f4 Qc7 8.Qf3 b5 9.Bxf6
B96.15=Sicilianskt: Najdorf, 7.f4 Nbd7
B96.16=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Bc4
B96.17=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qe2
B96.18=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qe2 Qc7
B96.19=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qf3
B96.20=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qf3 Qc7
B96.21=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qf3 Qc7 9.O-O-O b5
B96.22=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qf3 Qc7 9.O-O-O b5 10.Bd3
B96.23=Sicilianskt: Najdorf, 7.f4 Nbd7 8.Qf3 Qc7 9.O-O-O b5 10.e5
B96.24=Sicilianskt: Najdorf, Polugaevskyvarianten, 7.f4 b5
B96.25=Sicilianskt: Najdorf, Polugaevsky, 8.e5
B96.26=Sicilianskt: Najdorf, Polugaevsky, 9.fxe5 Qc7
B96.27=Sicilianskt: Najdorf, Polugaevsky, 10.Nf3
B96.28=Sicilianskt: Najdorf, Polugaevsky, 10.Bxb5+
B96.29=Sicilianskt: Najdorf, Polugaevsky, 10.exf6
B96.30=Sicilianskt: Najdorf, Polugaevsky, 10.exf6 Qe5+ 11.Be2
B96.31=Sicilianskt: Najdorf, Polugaevsky, 10.exf6 Qe5+ 11.Be2 Qxg5 12.Qd3
B96.32=Sicilianskt: Najdorf, Polugaevsky, 10.Qe2
B96.33=Sicilianskt: Najdorf, Polugaevsky, 10.Qe2 Nfd7 11.O-O-O Nc6
B96.34=Sicilianskt: Najdorf, Polugaevsky, 10.Qe2 Nfd7 11.O-O-O Bb7
B96.35=Sicilianskt: Najdorf, Polugaevsky, 10.Qe2 Nfd7 11.O-O-O Bb7 12.Qg4
B96.36=Sicilianskt: Najdorf, Polugaevsky, 10.Qe2 Nfd7 11.O-O-O Bb7 12.Qg4 Qxe5
B97.1=Sicilianskt: Najdorf, F�rgiftad bonde, 1.e4 c5 2.Nf3 d6 3.d4 cxd4 4.Nxd4 Nf6 5.Nc3 a6 6.Bg5 e6 7.f4 Qb6
B97.2=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Bxf6
B97.3=Sicilianskt: Najdorf, F�rgiftad bonde, 8.a3
B97.4=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Qd3
B97.5=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Nb3
B97.6=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Nb3 Be7
B97.7=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Nb3 Nbd7 9.Qf3
B97.8=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Nb3 Nbd7 9.Qf3 Be7
B97.9=Sicilianskt: Najdorf, F�rgiftad bonde, 8.Qd2
B97.10=Sicilianskt: Najdorf, Antagen F�rgiftad bonde, 8.Qd2 Qxb2
B97.11=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Nb3
B97.12=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Nb3 Nc6
B97.13=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Nb3 Qa3
B97.14=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Nb3 Qa3 10.Bxf6
B97.15=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Rb1
B97.16=Sicilianskt: Najdorf, F�rgiftad bonde, 9.Rb1 Qa3
B97.17=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Be2
B97.18=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Be2 Be7 11.O-O
B97.19=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Be2 Be7 11.O-O Nbd7
B97.20=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Bxf6
B97.21=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Bxf6 gxf6 11.Be2 Nc6
B97.22=Sicilianskt: Najdorf, F�rgiftad bonde, 10.Bxf6 gxf6 11.Be2 Bg7
B97.23=Sicilianskt: Najdorf, F�rgiftad bonde, 10.e5
B97.24=Sicilianskt: Najdorf, F�rgiftad bonde, 10.e5 dxe5
B97.25=Sicilianskt: Najdorf, F�rgiftad bonde, 10.e5 dxe5 11.fxe5 Nfd7 12.Bc4
B97.26=Sicilianskt: Najdorf, F�rgiftad bonde, 10.e5 dxe5 11.fxe5 Nfd7 12.Bc4 Bb4
B97.27=Sicilianskt: Najdorf, F�rgiftad bonde, 10.f5
B97.28=Sicilianskt: Najdorf, F�rgiftad bonde, 10.f5 Nc6
B97.29=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 7.f4 Qb6 8.Qd2 Qxb2 9.Rb1 Qa3 10.f5 Nc6 11.fxe6 fxe6 12.Nxc6 bxc6
B97.30=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, Timmans 13.Be2
B97.31=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5
B97.32=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 Nd5
B97.33=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5
B97.34=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5: 15.Ne4
B97.35=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5: 15.Ne4 Qxa2
B97.36=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5: 15.Ne4 Be7
B97.37=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5 med 18.c4
B97.38=Sicilianskt: Najdorf, F�rgiftad bonde, Huvudvarianten, 13.e5 dxe5 med 18.Nxf6+
B98.1=Sicilianskt: Najdorf, 7...Be7
B98.2=Sicilianskt: Najdorf, 7...Be7 8.Qf3
B98.3=Sicilianskt: Najdorf, Dannervarianten, 8.Qf3 Qa5
B98.4=Sicilianskt: Najdorf, Danner, 8.Qf3 Qa5 9.O-O-O Bd7
B98.5=Sicilianskt: Najdorf, Danner, 8.Qf3 Qa5 9.O-O-O Bd7 10.e5
B98.6=Sicilianskt: Najdorf, 7...Be7 8.Qf3 h6
B98.7=Sicilianskt: Najdorf, Brownevarianten, 8.Qf3 h6
B98.8=Sicilianskt: Najdorf, Browne, 10.O-O-O Nbd7
B98.9=Sicilianskt: Najdorf, Browne, 10.O-O-O Nbd7 11.Qg3
B98.10=Sicilianskt: Najdorf, Browne, 10.O-O-O Nbd7 11.Be2
B98.11=Sicilianskt: Najdorf, G�tenborg (Argentina)varianten, 8.Qf3 h6 9.Bh4 g5
B98.12=Sicilianskt: Najdorf, G�teborg, 11.Nxe6
B98.13=Sicilianskt: Najdorf, G�teborg, 11.Qh5
B98.14=Sicilianskt: Najdorf, 8...Qc7
B98.15=Sicilianskt: Najdorf, 8...Qc7 9.O-O-O Nc6
B99.1=Sicilianskt: Najdorf, Huvudvarianten, 8.Qf3 Qc7 9.O-O-O Nbd7
B99.2=Sicilianskt: Najdorf, Huvudvarianten, 10.Qg3
B99.3=Sicilianskt: Najdorf, Huvudvarianten, Keresvarianten, 10.Be2
B99.4=Sicilianskt: Najdorf, Huvudvarianten, Keres 10...b5 11.Bxf6 Nxf6 12.e5 Bb7
B99.5=Sicilianskt: Najdorf, Huvudvarianten, Keres, Queen Sacrifice Line, 10.Be2 b5 11.Bxf6 Nxf6 12.e5 Bb7 13.exf6
B99.6=Sicilianskt: Najdorf, Huvudvarianten, Keres, 13.Qg3
B99.7=Sicilianskt: Najdorf, Huvudvarianten, Keres, 13.Qg3 dxe5 14.fxe5 Nd7 15.Bxb5
B99.8=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3
B99.9=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 h6
B99.10=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 h6 11.Qh3
B99.11=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 h6 11.Bh4
B99.12=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 h6 11.Bh4 g5
B99.13=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 h6 11.Bh4 g5 12.fxg5
B99.14=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 b5
B99.15=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 b5 11.Rhe1 Bb7
B99.16=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 b5 11.Rhe1 Bb7 12.Nd5
B99.17=Sicilianskt: Najdorf, Huvudvarianten, 10.Bd3 b5 11.Rhe1 Bb7 12.Qg3
B99.18=Sicilianskt: Najdorf, Huvudvarianten, 10.g4
B99.19=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 h6
B99.20=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5
B99.21=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bd3
B99.22=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bd3 Bb7
B99.23=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.a3
B99.24=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bxf6
B99.25=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bxf6 gxf6
B99.26=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bxf6 Nxf6
B99.27=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bxf6 Nxf6 12.g5
B99.28=Sicilianskt: Najdorf, Huvudvarianten, 10.g4 b5 11.Bxf6 Nxf6 12.g5 Nd7 13.a3
B99.29=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5
B99.30=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5 Bxg5+
B99.31=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5 Bxg5+ 14.Kb1 Ne5
B99.32=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5 Nc5
B99.33=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5 Nc5 14.h4
B99.34=Sicilianskt: Najdorf, Moderna Huvudvarianten 13.f5 Nc5 14.f6
B99.35=Sicilianskt: Najdorf, Moderna Huvudvarianten, Perenyi, 13.f5 Nc5 14.f6 gxf6 15.gxf6 Bf8 16.Rg1
C00.1=Franskt:1.e4 e6
C00.2=Franskt:Birdvarianten, 1.e4 e6 2.Bb5
C00.3=Franskt:Reti (Spielmann)varianten, 1.e4 e6 2.b3
C00.4=Franskt:La Bourdonnaisvarianten, 1.e4 e6 2.f4
C00.5=Franskt:Steinitz attack, 1.e4 e6 2.e5
C00.6=Franskt:Steiner (Engelsk-Franska)varianten, 1.e4 e6 2.c4
C00.7=Franskt:Steiner (Engelsk-Franska)varianten, 1.e4 e6 2.c4 d5
C00.8=Franskt:Orthoschnapps gambit, 1.e4 e6 2.c4 d5 3.cxd5 exd5 4.Qb3
C00.9=Franskt:2.Nc3
C00.10=Franskt:2.Nc3 d5
C00.11=Franskt:Pelikanvarianten, 1.e4 e6 2.Nc3 d5 3.f4
C00.12=Franskt:Chigorinvarianten, 1.e4 e6 2.Qe2
C00.13=Franskt:Chigorin, 2...c5
C00.14=Franskt:Chigorin, 2...c5 3.Nf3
C00.15=Franskt:2.Nf3
C00.16=Franskt:2.Nf3 d5
C00.17=Franskt:2.Nf3 d5 3.e5
C00.18=Franskt:2.Nf3 d5 3.e5 c5
C00.19=Franskt:Vinggambit, 1.e4 e6 2.Nf3 d5 3.e5 c5 4.b4
C00.20=Franskt:Tv� springarvarianten, 1.e4 e6 2.Nf3 d5 3.Nc3
C00.21=Franskt:Antagen Kungsindisk 2.d3
C00.22=Franskt:Antagen Kungsindisk 2.d3 d5
C00.23=Franskt:Antagen Kungsindisk 2.d3 d5 3.Qe2
C00.24=Franskt:Antagen Kungsindisk 2.d3 d5 3.Qe2 Nf6
C00.25=Franskt:Antagen Kungsindisk 2.d3 d5 3.Nd2
C00.26=Franskt:Antagen Kungsindisk 2.d3 d5 3.Nd2 c5
C00.27=Franskt:Antagen Kungsindisk 2.d3 d5 3.Nd2 Nf6
C00.28=Franskt:Antagen Kungsindisk, Omv�nd Philidor 1.e4 e6 2.d3 d5 3.Nd2 Nf6 4.Ngf3
C00.29=Franskt:Antagen Kungsindisk, Omv�nd Philidor, 4...b6
C00.30=Franskt:Antagen Kungsindisk, Omv�nd Philidor, 4...Nc6
C00.31=Franskt:Antagen Kungsindisk, Omv�nd Philidor, 4...Nc6 5.c3
C00.32=Franskt:2.d4
C00.33=Franskt:St. George, 1.e4 e6 2.d4 a6
C00.34=Franskt:Franco-Benoni, 1.e4 e6 2.d4 c5
C00.35=Franskt:2.d4 d5
C00.36=Franskt:Alapin-Diemers gambit, 1.e4 e6 2.d4 d5 3.Be3
C00.37=Franskt:Schlechter, 1.e4 e6 2.d4 d5 3.Bd3
C01.1=Franskt:Avbyte, 1.e4 e6 2.d4 d5 3.exd5
C01.2=Franskt:Avbyte, 1.e4 e6 2.d4 d5 3.exd5 Qxd5
C01.3=Franskt:Avbyte, 1.e4 e6 2.d4 d5 3.exd5 exd5
C01.4=Franskt:Avbyte, 4.c4
C01.5=Franskt:Avbyte, 4.c4 c6
C01.6=Franskt:Avbyte, 4.c4 Nf6
C01.7=Franskt:Avbyte, 4.c4 Nf6 5.Nf3
C01.8=Franskt:Avbyte, 4.c4 Nf6 5.Nc3
C01.9=Franskt:Avbyte, 4.c4 Nf6 5.Nc3 c6
C01.10=Franskt:Avbyte, 4.c4 Nf6 5.Nc3 Bb4
C01.11=Franskt:Avbyte, 4.c4 Nf6 5.Nc3 Bb4 6.Nf3
C01.12=Franskt:Avbyte, 4.c4 Nf6 5.Nc3 Be7
C01.13=Franskt:Avbyte, 4.c4 Nf6 5.Nc3 Be7 6.Nf3
C01.14=Franskt:Avbyte, 4.Bf4
C01.15=Franskt:Avbyte, 4.Bd3
C01.16=Franskt:Avbyte, 4.Bd3 Nc6
C01.17=Franskt:Avbyte, 4.Bd3 Bd6
C01.18=Franskt:Avbyte, 4.Nf3
C01.19=Franskt:Avbyte, 4.Nf3 Nf6
C01.20=Franskt:Avbyte, 4.Nf3 Nf6 5.Bd3
C01.21=Franskt:Avbyte, 4.Nf3 Bd6
C01.22=Franskt:Avbyte, 4.Nf3 Bd6 5.Bd3
C01.23=Franskt:Avbyte, 4.Nf3 Bd6 5.Bd3 Nf6
C01.24=Franskt:Avbyte, 4.Nf3 Bd6 5.c4
C01.25=Franskt:Avbyte, 4.Nc3
C01.26=Franskt:Avbyte, 4.Nc3 Nf6
C01.27=Franskt:Avbyte, 4.Nc3 Nf6 5.Nf3
C01.28=Franskt:Avbyte, Svenoniusvarianten, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Nf6 5.Bg5
C01.29=Franskt:Avbyte, Bogoljubowvarianten, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Nf6 5.Bg5 Nc6
C01.30=Franskt:Avbyte Winawer, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Bb4
C01.31=Franskt:Avbyte Winawer, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Bb4 5.Bd3
C01.32=Franskt:Avbyte, Canal attack, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Bb4 5.Bd3 Ne7 6.Qh5
C01.33=Franskt:Avbyte Winawer, 1.e4 e6 2.d4 d5 3.exd5 exd5 4.Nc3 Bb4 5.Bd3 Nc6
C02.1=Franskt:Avancera, 1.e4 e6 2.d4 d5 3.e5
C02.2=Franskt:Avancera, 3...Ne7
C02.3=Franskt:Avancera, 3...b6
C02.4=Franskt:Avancera, 3...b6
C02.5=Franskt:Avancera, 3...c5
C02.6=Franskt:Avancera, Vinggambit, 1.e4 e6 2.d4 d5 3.e5 c5 4.b4
C02.7=Franskt:Avancera, Steinitz, 1.e4 e6 2.d4 d5 3.e5 c5 4.dxc5
C02.8=Franskt:Avancera, Nimzowitschs attack, 1.e4 e6 2.d4 d5 3.e5 c5 4.Qg4
C02.9=Franskt:Avancera, Nimzowitschs gambit, 1.e4 e6 2.d4 d5 3.e5 c5 4.Qg4 cxd4 5.Nf3
C02.10=Franskt:Avancera, 4.Nf3
C02.11=Franskt:Avancera, Ruisdonks gambit, 1.e4 e6 2.d4 d5 3.e5 c5 4.Nf3 cxd4 5.Bd3
C02.12=Franskt:Avancera, 4.c3
C02.13=Franskt:Avancera, 4.c3 Qb6
C02.14=Franskt:Avancera, Wade, 1.e4 e6 2.d4 d5 3.e5 c5 4.c3 Qb6 5.Nf3 Bd7
C02.15=Franskt:Avancera, Wade, 6.Be2
C02.16=Franskt:Avancera, 4...Nc6
C02.17=Franskt:Avancera, Paulsen, 1.e4 e6 2.d4 d5 3.e5 c5 4.c3 Nc6 5.Nf3
C02.18=Franskt:Avancera, 5.Nf3 Nge7
C02.19=Franskt:Avancera, Euwe, 1.e4 e6 2.d4 d5 3.e5 c5 4.c3 Nc6 5.Nf3 Bd7
C02.20=Franskt:Avancera, Euwe, 6.a3
C02.21=Franskt:Avancera, Euwe, 6.Be2
C02.22=Franskt:Avancera, Euwe, 6.Be2 Nge7
C02.23=Franskt:Avancera, 5.Nf3 Qb6
C02.24=Franskt:Avancera, Milner-Barrys gambit, 1.e4 e6 2.d4 d5 3.e5 c5 4.c3 Nc6 5.Nf3 Qb6 6.Bd3
C02.25=Franskt:Avancera, 5.Nf3 Qb6 6.Be2
C02.26=Franskt:Avancera, 5.Nf3 Qb6 6.Be2 cxd4 7.cxd4
C02.27=Franskt:Avancera, 5.Nf3 Qb6 6.a3
C02.28=Franskt:Avancera, 5.Nf3 Qb6 6.a3 Bd7
C02.29=Franskt:Avancera, 5.Nf3 Qb6 6.a3 Nh6
C02.30=Franskt:Avancera, 5.Nf3 Qb6 6.a3 c4
C02.31=Franskt:Avancera, 5.Nf3 Qb6 6.a3 c4 7.Nbd2
C03.1=Franskt:Tarrasch, 1.e4 e6 2.d4 d5 3.Nd2
C03.2=Franskt:Tarrasch, 3...dxe4
C03.3=Franskt:Tarrasch, Haberditzvarianten, 1.e4 e6 2.d4 d5 3.Nd2 f5
C03.4=Franskt:Tarrasch, 3...b6
C03.5=Franskt:Tarrasch, 3...a6
C03.6=Franskt:Tarrasch, 3...a6 4.Ngf3
C03.7=Franskt:Tarrasch, 3...Be7
C03.8=Franskt:Tarrasch, 3...Be7 4.Bd3
C03.9=Franskt:Tarrasch, 3...Be7 4.Bd3 c5
C03.10=Franskt:Tarrasch, 3...Be7 4.Bd3 c5 5.dxc5 Nf6
C03.11=Franskt:Tarrasch, 3...Be7 4.Ngf3
C03.12=Franskt:Tarrasch, 3...Be7 4.Ngf3 Nf6
C03.13=Franskt:Tarrasch, 3...Be7 4.Ngf3 Nf6 5.Bd3
C03.14=Franskt:Tarrasch, Guimardvarianten, 1.e4 e6 2.d4 d5 3.Nd2 Nc6
C03.15=Franskt:Tarrasch, Guimard, 1.e4 e6 2.d4 d5 3.Nd2 Nc6 4.c3
C03.16=Franskt:Tarrasch, Guimard, 1.e4 e6 2.d4 d5 3.Nd2 Nc6 4.c3 e5
C03.17=Franskt:Tarrasch, Guimard, 1.e4 e6 2.d4 d5 3.Nd2 Nc6 4.Ngf3
C04.1=Franskt:Tarrasch, Guimard, 4.Ngf3 Nf6
C04.2=Franskt:Tarrasch, Guimard, 4.Ngf3 Nf6 5.e5
C04.3=Franskt:Tarrasch, Guimard, Huvudvarianten
C04.4=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.c3
C04.5=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Bb5
C04.6=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Be2
C04.7=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Be2 f6
C04.8=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Nb3
C04.9=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Nb3 a5
C04.10=Franskt:Tarrasch, Guimard, Huvudvarianten, 6.Nb3 Be7
C05.1=Franskt:Tarrasch, St�ngd, 1.e4 e6 2.d4 d5 3.Nd2 Nf6
C05.2=Franskt:Tarrasch, St�ngd, 4.e5
C05.3=Franskt:Tarrasch, St�ngd, 4...Ne4
C05.4=Franskt:Tarrasch, St�ngd, 4...Ne4 5.Nxe4
C05.5=Franskt:Tarrasch, St�ngd, 4...Nfd7
C05.6=Franskt:Tarrasch, St�ngd, 5.f4
C05.7=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6
C05.8=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3
C05.9=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 cxd4
C05.10=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6
C05.11=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.h4
C05.12=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.h4
C05.13=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.Ne2
C05.14=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.Ne2
C05.15=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.g3
C05.16=Franskt:Tarrasch, St�ngd, 5.f4 c5 6.c3 Nc6 7.Ndf3 Qb6 8.g3
C05.17=Franskt:Tarrasch, St�ngd, 5.c3
C05.18=Franskt:Tarrasch, 5.Bd3
C05.19=Franskt:Tarrasch, Botvinnik, 1.e4 e6 2.d4 d5 3.Nd2 Nf6 4.e5 Nfd7 5.Bd3 c5 6.c3 b6
C05.20=Franskt:Tarrasch, St�ngd, 6...Nc6
C05.21=Franskt:Tarrasch, St�ngd, 7.Ndf3
C05.22=Franskt:Tarrasch, St�ngd, 7.Ndf3 Qa5
C05.23=Franskt:Tarrasch, St�ngd, 7.Ngf3
C05.24=Franskt:Tarrasch, St�ngd, 7.Ngf3 Be7
C05.25=Franskt:Tarrasch, St�ngd, 7.Ngf3 Be7 8.O-O g5
C05.26=Franskt:Tarrasch, St�ngd, Nunn-Korchnois gambit, 4.e5 Nfd7 5.Bd3 c5 6.c3 Nc6 7.Ngf3 Qb6 8.O-O
C05.27=Franskt:Tarrasch, St�ngd, 7.Ne2
C05.28=Franskt:Tarrasch, St�ngd, 7.Ne2 a5
C06.1=Franskt:Tarrasch, St�ngd, Huvudvarianten, 3.Nd2 Nf6 4.e5 Nfd7 5.Bd3 c5 6.c3 Nc6 7.Ne2 cxd4 8.cxd4
C06.2=Franskt:Tarrasch, St�ngd, Leningrad, 3.Nd2 Nf6 4.e5 Nfd7 5.Bd3 c5 6.c3 Nc6 7.Ne2 cxd4 8.cxd4 Nb6
C06.3=Franskt:Tarrasch, St�ngd, Leningrad, 9.Nf3
C06.4=Franskt:Tarrasch, St�ngd, Leningrad, 9.O-O
C06.5=Franskt:Tarrasch, St�ngd, Leningrad, 9.O-O a5
C06.6=Franskt:Tarrasch, St�ngd, Leningrad, 9.O-O Bd7
C06.7=Franskt:Tarrasch, St�ngd, 8...Qb6
C06.8=Franskt:Tarrasch, St�ngd, 8...Qb6 9.O-O
C06.9=Franskt:Tarrasch, St�ngd, 8...Qb6 9.Nf3
C06.10=Franskt:Tarrasch, St�ngd, 8...Qb6 9.Nf3 f6
C06.11=Franskt:Tarrasch, St�ngd, 8...f6
C06.12=Franskt:Tarrasch, St�ngd, 8...f6 9.Nf4
C06.13=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6
C06.14=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6 Nxf6
C06.15=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6 Nxf6 10.O-O Bd6 11.Nf3
C06.16=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...Qb6
C06.17=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...Qb6 12.Nc3
C06.18=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...Qc7
C06.19=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...Qc7 12.Bg5
C06.20=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...O-O
C06.21=Franskt:Tarrasch, St�ngd, 8...f6 9.exf6, 11...O-O 12.Bf4
C07.1=Franskt:Tarrasch, �ppen, 1.e4 e6 2.d4 d5 3.Nd2 c5
C07.2=Franskt:Tarrasch, �ppen, 4.c3
C07.3=Franskt:Tarrasch, �ppen, 4.dxc5
C07.4=Franskt:Tarrasch, �ppen, 4.Ngf3
C07.5=Franskt:Tarrasch, �ppen, 4.Ngf3 a6
C07.6=Franskt:Tarrasch, �ppen, 4.Ngf3 Nf6
C07.7=Franskt:Tarrasch, �ppen, 4.Ngf3 Nc6
C07.8=Franskt:Tarrasch, �ppen, 4.Ngf3 cxd4
C07.9=Franskt:Tarrasch, �ppen, 4.exd5
C07.10=Franskt:Tarrasch, Shaposhnikovs gambit, 1.e4 e6 2.d4 d5 3.Nd2 c5 4.exd5 Nf6
C07.11=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5
C07.12=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5 5.Ngf3
C07.13=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5 5.Ngf3 cxd4
C07.14=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5 5.Ngf3 cxd4 6.Bc4
C07.15=Franskt:Tarrasch, �ppen, Eliskasesvarianten, 1.e4 e6 2.d4 d5 3.Nd2 c5 4.exd5 Qxd5 5.Ngf3 cxd4 6.Bc4 Qd8
C07.16=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5 5.Ngf3 cxd4 6.Bc4 Qd6
C07.17=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Qxd4
C07.18=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Qxd4 Qxd4
C07.19=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Nxd4
C07.20=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Nxd4 a6
C07.21=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Nxd4 a6 11.c3
C07.22=Franskt:Tarrasch, �ppen, 4.exd5 Qxd5, Huvudvarianten, 10.Nxd4 a6 11.Re1
C08.1=Franskt:Tarrasch, �ppen, 4.exd5 exd5
C08.2=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Bb5+ Nc6
C08.3=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Bb5+ Nc6 6.Qe2+
C08.4=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Bb5+ Bd7
C08.5=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Bb5+ Bd7 6.Qe2+
C08.6=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Bb5+ Bd7 6.Qe2+ Be7
C08.7=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Ngf3
C08.8=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Ngf3 a6
C08.9=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Ngf3 a6 6.Be2
C08.10=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Ngf3 Nf6
C08.11=Franskt:Tarrasch, �ppen, 4.exd5 exd5 5.Ngf3 Nf6, 7.Bxd7
C08.12=Franskt:Tarrasch, �ppen, Huvudvarianten, 4.exd5 exd5 5.Ngf3 Nf6
C08.13=Franskt:Tarrasch, �ppen, Huvudvarianten, 4.exd5 exd5 5.Ngf3 Nf6, 10.Nb3
C09.1=Franskt:Tarrasch, �ppen, 5.Ngf3 Nc6
C09.2=Franskt:Tarrasch, �ppen, 5.Ngf3 Nc6 6.Bb5
C09.3=Franskt:Tarrasch, �ppen, 5.Ngf3 Nc6 6.Bb5 cxd4
C09.4=Franskt:Tarrasch, �ppen, 5.Ngf3 Nc6 6.Bb5 Bd6
C09.5=Franskt:Tarrasch, �ppen, 7.O-O
C09.6=Franskt:Tarrasch, �ppen, 7.dxc5
C09.7=Franskt:Tarrasch, �ppen, Huvudvarianten, 6.Bb5 Bd6 7.dxc5 Bxc5 8.O-O Ne7
C09.8=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.c3
C09.9=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.c3 O-O 10.Nb3 Bd6
C09.10=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.c3 O-O 10.Nb3 Bb6
C09.11=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.c3 O-O 10.Nb3 Bb6 11.Re1
C09.12=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3
C09.13=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bb6
C09.14=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6
C09.15=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6 10.Nbd4
C09.16=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6 10.Bg5
C09.17=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6 10.Re1
C09.18=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6 10.Re1 O-O 11.Bg5
C09.19=Franskt:Tarrasch, �ppen, Huvudvarianten, 9.Nb3 Bd6 10.Re1 O-O 11.Bg5 Bg4
C10.1=Franskt:1.e4 e6 2.d4 d5 3.Nc3
C10.2=Franskt:Marshallvarianten, 1.e4 e6 2.d4 d5 3.Nc3 c5
C10.3=Franskt:3.Nc3 Nc6
C10.4=Franskt:3.Nc3 Nc6 4.Nf3 Nf6
C10.5=Franskt:3.Nc3 Be7
C10.6=Franskt:Rubinstein, 1.e4 e6 2.d4 d5 3.Nc3 dxe4
C10.7=Franskt:Rubinstein, 1.e4 e6 2.d4 d5 3.Nc3 dxe4 4.Nxe4
C10.8=Franskt:Rubinstein, Ellis gambit, 1.e4 e6 2.d4 d5 3.Nc3 dxe4 4.Nxe4 e5
C10.9=Franskt:Rubinstein, Frere (Becker)varianten, 1.e4 e6 2.d4 d5 3.Nc3 dxe4 4.Nxe4 Qd5
C10.10=Franskt:Rubinstein, 4...Nf6
C10.11=Franskt:Rubinstein, 4...Nd7
C10.12=Franskt:Rubinstein, 5.Nf3 Be7
C10.13=Franskt:Rubinstein, 5.Nf3 Ngf6
C10.14=Franskt:Rubinstein, 5.Nf3 Ngf6 6.Bd3
C10.15=Franskt:Rubinstein, 5.Nf3 Ngf6 6.Nxf6+
C10.16=Franskt:Rubinstein, Capablanca, 3.Nc3 dxe4 4.Nxe4 Nd7 5.Nf3 Ngf6 6.Nxf6+ Nxf6 7.Ne5
C10.17=Franskt:Rubinstein, 7.Bd3
C10.18=Franskt:Rubinstein, 7.Bd3 c5
C10.19=Franskt:Rubinstein, 7.Bd3 c5 8.dxc5
C10.20=Franskt:Rubinstein, 7.Bg5
C10.21=Franskt:Rubinstein, 4...Bd7
C10.22=Franskt:Rubinstein, 4...Bd7 5.Nf3
C10.23=Franskt:Rubinstein, 4...Bd7 5.Nf3 Bc6 6.Bd3
C10.24=Franskt:Rubinstein, 4...Bd7 5.Nf3 Bc6 6.Bd3 Nd7
C10.25=Franskt:Rubinstein, 4...Bd7 5.Nf3 Bc6 6.Bd3 Nd7 7.O-O
C10.26=Franskt:Rubinstein, 4...Bd7 5.Nf3 Bc6 6.Bd3 Nd7 7.O-O Ngf6
C10.27=Franskt:Rubinstein, 4...Bd7 5.Nf3 Bc6 6.Bd3 Nd7 7.O-O Ngf6 8.Ng3
C11.1=Franskt:3.Nc3 Nf6
C11.2=Franskt:Hennebergervarianten, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.Be3
C11.3=Franskt:3.Nc3 Nf6 4.exd5
C11.4=Franskt:Schweiziskvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.Bd3
C11.5=Franskt:Steinitz
C11.6=Franskt:Steinitz, Gledhill attack, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.e5 Nfd7 5.Qg4
C11.7=Franskt:Steinitz, 5.Nf3
C11.8=Franskt:Steinitz, 5.Nf3 c5
C11.9=Franskt:Steinitz, 5.Nf3 c5 6.dxc5
C11.10=Franskt:Steinitz, 5.f4
C11.11=Franskt:Steinitz, 5.f4 c5
C11.12=Franskt:Steinitz, 6.dxc5
C11.13=Franskt:Steinitz, Bradford attack, 4.e5 Nfd7 5.f4 c5 6.dxc5 Bxc5 7.Qg4
C11.14=Franskt:Steinitz, 6.dxc5 Nc6
C11.15=Franskt:Steinitz, Brodsky-Jonesvarianten, 4.e5 Nfd7 5.f4 c5 6.dxc5 Nc6 7.a3 Bxc5 8.Qg4 O-O 9.Nf3 f6
C11.16=Franskt:Steinitz, 6.Nf3
C11.17=Franskt:Steinitz, BoleSlaviskskyvarianten, 4.e5 Nfd7 5.f4 c5 6.Nf3 Nc6 7.Be3
C11.18=Franskt:Steinitz, BoleSlavisksky, 7...a6
C11.19=Franskt:Steinitz, BoleSlavisksky, 7...a6 8.Qd2 b5
C11.20=Franskt:Steinitz, BoleSlavisksky, 7...cxd4
C11.21=Franskt:Steinitz, BoleSlavisksky, 7...cxd4 8.Nxd4 Qb6
C11.22=Franskt:Steinitz, BoleSlavisksky, 7...cxd4 8.Nxd4 Bc5
C11.23=Franskt:3.Nc3 Nf6 4.Bg5
C11.24=Franskt:Burnvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.Bg5 dxe4
C11.25=Franskt:Burn, 5.Nxe4
C11.26=Franskt:Burn, 5.Nxe4 Nbd7
C11.27=Franskt:Burn, 5.Nxe4 Nbd7 6.Nf3
C11.28=Franskt:Burn, 5.Nxe4 Nbd7 6.Nf3 Be7
C11.30=Franskt:Burn, 5.Nxe4 Be7
C11.31=Franskt:Burn, 6.Bxf6 Bxf6
C11.32=Franskt:Burn, 6.Bxf6 gxf6
C11.33=Franskt:Burn, 6.Bxf6 gxf6 7.Nf3
C11.34=Franskt:Burn, 6.Bxf6 gxf6 7.Nf3 b6
C11.35=Franskt:Burn, 6.Bxf6 gxf6 7.Nf3 b6 8.Bd3
C11.36=Franskt:Burn, 6.Bxf6 gxf6 7.Nf3 b6 8.Bc4
C11.37=Franskt:Burn, 6.Bxf6 gxf6 7.Nf3 f5
C12.1=Franskt:MacCutcheon, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.Bg5 Bb4
C12.2=Franskt:MacCutcheon, 5.exd5
C12.3=Franskt:MacCutcheon, 5.exd5 Qxd5
C12.4=Franskt:MacCutcheon, Bogoljubowvarianten, 5.exd5 Qxd5 6.Bxf6 gxf6 7.Qd2 Qa5
C12.5=Franskt:MacCutcheon, Avanceravarianten, 5.e5
C12.6=Franskt:MacCutcheon, Avanceravarianten, 5.e5 h6
C12.7=Franskt:MacCutcheon, Chigorinvarianten, 5.e5 h6 6.exf6
C12.8=Franskt:MacCutcheon, Grigorievvarianten, 5.e5 h6 6.exf6 hxg5 7.fxg7 Rg8 8.h4 gxh4 9.Qg4
C12.9=Franskt:MacCutcheon, Olland (Holl�ndsk)varianten, 5.e5 h6 6.Bc1
C12.10=Franskt:MacCutcheon, Bernsteinvarianten, 5.e5 h6 6.Bh4
C12.11=Franskt:MacCutcheon, Janowskivarianten, 5.e5 h6 6.Be3
C12.12=Franskt:MacCutcheon, 6.Bd2
C12.13=Franskt:MacCutcheon, Tartakowervarianten, 5.e5 h6 6.Bd2 Nfd7
C12.14=Franskt:MacCutcheon, Laskervarianten, 5.e5 h6 6.Bd2 Bxc3
C12.15=Franskt:MacCutcheon, Lasker, 7.bxc3
C12.16=Franskt:MacCutcheon, 8.Qg4
C12.17=Franskt:MacCutcheon, 8.Qg4 Kf8
C12.18=Franskt:MacCutcheon, Durasvarianten, 5.e5 h6 6.Bd2 Bxc3 7.bxc3 Ne4 8.Qg4 Kf8 9.Bc1
C12.19=Franskt:MacCutcheon, 8.Qg4 Kf8 9.Bd3
C12.20=Franskt:MacCutcheon, 8.Qg4 g6
C12.21=Franskt:MacCutcheon, 8.Qg4 g6 9.Bd3
C12.22=Franskt:MacCutcheon, Huvudvarianten, 5.e5 h6 6.Bd2 Bxc3 7.bxc3 Ne4 8.Qg4 g6 9.Bd3 Nxd2 10.Kxd2 c5
C12.23=Franskt:MacCutcheon, Huvudvarianten, 11.Nf3
C12.24=Franskt:MacCutcheon, Huvudvarianten, 11.Nf3 Nc6
C13.1=Franskt:Klassisk, 1.e4 e6 2.d4 d5 3.Nc3 Nf6 4.Bg5 Be7
C13.2=Franskt:Klassisk, Anderssenvarianten, 5.Bxf6
C13.3=Franskt:Klassisk, Anderssen-Richtervarianten, 5.Bxf6 Bxf6 6.e5 Be7 7.Qg4
C13.4=Franskt:Klassisk, 5.e5
C13.5=Franskt:Klassisk, Nimzowitschvarianten, 5.e5 Ng8
C13.6=Franskt:Klassisk, Frankfurtvarianten, 5.e5 Ng8 6.Be3 b6
C13.7=Franskt:Klassisk, Tartakowervarianten, 5.e5 Ne4
C13.8=Franskt:Klassisk, Tartakower, 6.Bxe7
C13.9=Franskt:Klassisk, 5.e5 Nfd7
C13.10=Franskt:Chatard-Alekhine attack, 5.e5 Nfd7
C13.11=Franskt:Chatard-Alekhine, Teichmannvarianten, 5.e5 Nfd7 6.h4 f6
C13.12=Franskt:Chatard-Alekhine, Spielmannvarianten, 5.e5 Nfd7 6.h4 O-O
C13.13=Franskt:Chatard-Alekhine, 6...Bxg5
C13.14=Franskt:Chatard-Alekhine, 6...Bxg5 7.hxg5 Qxg5
C13.15=Franskt:Chatard-Alekhine, 6...Bxg5 7.hxg5 Qxg5 8.Nh3 Qe7 9.Nf4
C13.16=Franskt:Chatard-Alekhine, Maroczyvarianten, 5.e5 Nfd7 6.h4 a6
C13.17=Franskt:Chatard-Alekhine, Maroczy, 7.Qg4 Bxg5
C13.18=Franskt:Chatard-Alekhine, Breyervarianten, 5.e5 Nfd7 6.h4 c5
C13.19=Franskt:Chatard-Alekhine, Breyer, 7.Bxe7
C13.20=Franskt:Chatard-Alekhine, Breyer, 7.Bxe7 Kxe7
C14.1=Franskt:Klassisk, 6.Bxe7 Qxe7
C14.2=Franskt:Klassisk, Pollockvarianten, 7.Qg4
C14.3=Franskt:Klassisk, Tarraschvarianten, 7.Bd3
C14.4=Franskt:Klassisk, Alapinvarianten, 7.Nb5
C14.5=Franskt:Klassisk, Rubinsteinvarianten, 7.Qd2
C14.6=Franskt:Klassisk, Steinitzvarianten, 7.f4
C14.7=Franskt:Klassisk, Steinitz, 7...a6
C14.8=Franskt:Klassisk, Steinitz, 7...a6 8.Nf3 c5
C14.9=Franskt:Klassisk, Steinitz, 7...a6 8.Nf3 c5
C14.10=Franskt:Klassisk, Steinitz, 7...O-O
C14.11=Franskt:Klassisk, Steinitz, 7...O-O 8.Nf3 c5
C14.12=Franskt:Klassisk, Steinitz, 8.Nf3 c5 9.dxc5
C14.13=Franskt:Klassisk, Steinitz, 9.Qd2
C14.14=Franskt:Klassisk, St�hlbergvarianten, 7.f4 O-O 8.Nf3 c5 9.Qd2 Nc6 10.O-O-O c4
C14.15=Franskt:Klassisk, Steinitz, 9.Qd2 Nc6 10.dxc5
C14.16=Franskt:Klassisk, Steinitz, 9.Qd2 Nc6 10.dxc5 Qxc5
C15.1=Franskt:Winawer, 1.e4 e6 2.d4 d5 3.Nc3 Bb4
C15.2=Franskt:Winawer, 4.exd5
C15.4=Franskt:Winawer, 4.Qg4
C15.5=Franskt:Winawer, 4.Qd3
C15.6=Franskt:Winawer, 4.Qd3 dxe4
C15.7=Franskt:Winawer, 4.Bd3
C15.8=Franskt:Winawer, 4.Bd3 c5
C15.9=Franskt:Winawer, Kondratiyevvarianten, 4.Bd3 c5 5.exd5 Qxd5 6.Bd2
C15.10=Franskt:Winawer, 4.Bd3 dxe4
C15.11=Franskt:Winawer, 4.Bd3 dxe4 5.Bxe4
C15.12=Franskt:Winawer, 4.Bd3 dxe4 5.Bxe4 Nf6
C15.13=Franskt:Winawer, M�ller-Zhuravlevs gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.Bd2
C15.14=Franskt:Winawer, M�ller-Zhuravlevs gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.Bd2 dxe4
C15.15=Franskt:Winawer, M�ller-Zhuravlevs gambit, 5.Qg4
C15.16=Franskt:Winawer, M�ller-Zhuravlevs gambit, Kuninvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.Bd2 dxe4 5.Qg4 Qxd4
C15.17=Franskt:Winawer, M�ller-Zhuravlevs gambit, 5.Qg4 Nf6
C15.18=Franskt:Winawer, 4.a3
C15.19=Franskt:Winawer, 4.a3 Bxc3+
C15.20=Franskt:Winawer, 4.a3 Bxc3+
C15.21=Franskt:Winawer, 4.a3 Bxc3+ 5.bxc3 dxe4
C15.22=Franskt:Winawer, Winkelmann-Reimers gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.a3 Bxc3+ 5.bxc3 dxe4 6.f3
C15.23=Franskt:Winawer, Antagen Winkelmann-Reimers gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.a3 Bxc3+ 5.bxc3 dxe4 6.f3 exf3
C15.24=Franskt:Winawer, Winkelmann-Reimer, H�bner f�rsvar, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.a3 Bxc3+ 5.bxc3 dxe4 6.f3 e5
C15.25=Franskt:Winawer, Winkelmann-Reimer, 6...c5
C15.26=Franskt:Winawer, 4.a3 Bxc3+ 5.bxc3 dxe4 6.Qg4
C15.27=Franskt:Winawer, Alekhines gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.Ne2
C15.28=Franskt:Winawer, Alekhines gambit, 4...Nf6
C15.29=Franskt:Winawer, Alekhines gambit, 4...Nc6
C15.30=Franskt:Winawer, Antagen Alekhines gambit, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.Ne2 dxe4
C15.31=Franskt:Winawer, Alekhines gambit, 5.a3 Bxc3+
C15.32=Franskt:Winawer, Alekhines gambit, Kanvarianten
C15.33=Franskt:Winawer, Alekhines gambit, Kan, 7.Bb5
C15.34=Franskt:Winawer, Alekhines gambit, 5.a3 Be7
C15.35=Franskt:Winawer, Alekhines gambit, 5.a3 Be7 6.Nxe4 Nf6
C15.36=Franskt:Winawer, Alekhines gambit, Alatortsevvarianten, 4.Ne2 dxe4 5.a3 Be7 6.Nxe4 Nf6 7.N2g3 O-O 8.Be2 Nc6
C15.37=Franskt:Winawer, Alekhines gambit, 5.a3 Be7 6.Nxe4 Nf6 7.Qd3
C16.1=Franskt:Winawer, Avanceravarianten, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.e5
C16.2=Franskt:Winawer, 4.e5 b6
C16.3=Franskt:Winawer, 4.e5 b6 5.Qg4
C16.4=Franskt:Winawer, 4.e5 b6 5.Qg4 Bf8 6.Bg5
C16.5=Franskt:Winawer, 4.e5 b6 5.a3
C16.6=Franskt:Winawer, 4.e5 b6 5.a3 Bf8
C16.7=Franskt:Winawer, Petrosianvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.e5 Qd7
C16.8=Franskt:Winawer, Petrosian, 5.Bd2
C16.9=Franskt:Winawer, Petrosian, 5.a3
C16.10=Franskt:Winawer, Petrosian, 5.a3 Bxc3+ 6.bxc3 b6
C16.11=Franskt:Winawer, Petrosian, 5.a3 Bxc3+ 6.bxc3 b6 7.Qg4
C16.12=Franskt:Winawer, Avancera, 4...Ne7
C16.13=Franskt:Winawer, Avancera, 4...Ne7 5.Bd2
C16.14=Franskt:Winawer, Avancera, 4...Ne7 5.Bd2 b6
C16.15=Franskt:Winawer, Avancera, 4...Ne7 5.a3
C16.16=Franskt:Winawer, Avancera, 4...Ne7 5.a3 Bxc3+ 6.bxc3 b6
C16.17=Franskt:Winawer, Avancera, 4...Ne7 5.a3 Bxc3+ 6.bxc3 b6 7.Qg4
C17.1=Franskt:Winawer, Avancera, 4...c5
C17.2=Franskt:Winawer, Avancera, 5.dxc5
C17.3=Franskt:Winawer, Ryska varianten, 5.Qg4
C17.4=Franskt:Winawer, Rysk, 5.Qg4 Ne7 6.dxc5
C17.5=Franskt:Winawer, Bogoljubowvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.e5 c5 5.Bd2
C17.6=Franskt:Winawer, Bogoljubow, 5...cxd4
C17.7=Franskt:Winawer, Bogoljubow, 5...Ne7
C17.8=Franskt:Winawer, Bogoljubow, 5...Ne7 6.a3
C17.9=Franskt:Winawer, Bogoljubow, 5...Ne7 6.dxc5
C17.10=Franskt:Winawer, Bogoljubow, 5...Ne7 6.Nb5
C17.11=Franskt:Winawer, 5.a3
C17.12=Franskt:Winawer, 5.a3 cxd4
C17.13=Franskt:Winawer, Rauzervarianten, 5.a3 cxd4 6.axb4 dxc3 7.Nf3
C17.14=Franskt:Winawer, Schweiziska varianten, 5.a3 Ba5
C17.15=Franskt:Winawer, Schweizisk, 6.b4
C17.16=Franskt:Winawer, Schweizisk, 6.b4 cxd4 7.Qg4
C17.17=Franskt:Winawer, Schweizisk, 6.b4 cxd4 7.Qg4 Ne7 8.bxa5
C17.18=Franskt:Winawer, Schweizisk, 6.b4 cxd4 7.Nb5
C17.19=Franskt:Winawer, Schweizisk, 6.b4 cxd4 7.Nb5 Bc7 8.f4
C17.20=Franskt:Winawer, Schweizisk, 6.b4 cxd4 7.Nb5 Bc7 8.f4 Bd7
C18.1=Franskt:Winawer, 5...Bxc3+
C18.2=Franskt:Winawer, 5...Bxc3+ 6.bxc3
C18.3=Franskt:Winawer, 6...Qa5
C18.4=Franskt:Winawer, 6...Qc7
C18.5=Franskt:Winawer, 6...Qc7 7.Qg4
C18.6=Franskt:Winawer, 6...Qc7 7.Qg4 f6
C18.7=Franskt:Winawer, 6...Qc7 7.Qg4 f5
C18.8=Franskt:Winawer, 6...Ne7
C18.9=Franskt:Winawer, 6...Ne7 7.h4
C18.10=Franskt:Winawer, 6...Ne7 7.h4 Qc7
C18.12=Franskt:Winawer, 6...Ne7 7.h4 Nbc6
C18.13=Franskt:Winawer, 6...Ne7 7.h4 Nbc6 8.Nf3
C18.14=Franskt:Winawer, 6...Ne7 7.Qg4
C18.15=Franskt:Winawer, 6...Ne7 7.Qg4 Nbc6
C18.16=Franskt:Winawer, 6...Ne7 7.Qg4 Kf8
C18.17=Franskt:Winawer, 6...Ne7 7.Qg4 cxd4
C18.18=Franskt:Winawer, 6...Ne7 7.Qg4 O-O
C18.19=Franskt:Winawer, 6...Ne7 7.Qg4 O-O 8.Bd3
C18.20=Franskt:Winawer, 6...Ne7 7.Qg4 O-O 8.Bd3 Nbc6
C18.21=Franskt:Winawer, 6...Ne7 7.Qg4 O-O 8.Nf3
C18.22=Franskt:Winawer, 6...Ne7 7.Qg4 O-O 8.Nf3 Nbc6
C18.23=Franskt:Winawer, F�rgiftad bonde, 6.bxc3 Ne7 7.Qg4 Qc7
C18.24=Franskt:Winawer, F�rgiftad bonde, 8.Qxg7
C18.25=Franskt:Winawer, F�rgiftad bonde, 10.Qd3
C18.26=Franskt:Winawer, F�rgiftad bonde, Euwe-Gligoricvarianten, 6.bxc3 Ne7 7.Qg4 Qc7 8.Qxg7 Rg8 9.Qxh7 cxd4 10.Kd1
C18.27=Franskt:Winawer, F�rgiftad bonde, Konstantinopolskyvarianten, 6.bxc3 Ne7 7.Qg4 Qc7 8.Qxg7 Rg8 9.Qxh7 cxd4 10.Ne2
C18.28=Franskt:Winawer, F�rgiftad bonde, Huvudvarianten, 10.Ne2 Nbc6 11.f4 Bd7 12.Qd3 dxc3
C18.29=Franskt:Winawer, F�rgiftad bonde, Huvudvarianten, 13.Nxc3
C19.1=Franskt:Winawer, Smyslovvarianten, 1.e4 e6 2.d4 d5 3.Nc3 Bb4 4.e5 c5 5.a3 Bxc3+ 6.bxc3 Ne7 7.a4
C19.2=Franskt:Winawer, Smyslov, 7...Qa5
C19.3=Franskt:Winawer, 6...Ne7 7.Nf3
C19.4=Franskt:Winawer, 6...Ne7 7.Nf3 Qc7
C19.5=Franskt:Winawer, 6...Ne7 7.Nf3 Qc7 8.a4
C19.6=Franskt:Winawer, 6...Ne7 7.Nf3 Qc7 8.a4 b6
C19.7=Franskt:Winawer, 6...Ne7 7.Nf3 Qa5
C19.8=Franskt:Winawer, 6...Ne7 7.Nf3 b6
C19.9=Franskt:Winawer, 6...Ne7 7.Nf3 b6 8.a4
C19.10=Franskt:Winawer, 6...Ne7 7.Nf3 b6 8.Bb5+
C19.11=Franskt:Winawer, 6...Ne7 7.Nf3 Bd7
C19.12=Franskt:Winawer, 6...Ne7 7.Nf3 Bd7 8.a4
C19.13=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6
C19.14=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4
C19.15=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Bd7
C19.16=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5
C19.17=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5 9.Qd2
C19.18=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5 9.Qd2 Bd7
C19.19=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5+ 9.Bd2
C19.20=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5+ 9.Bd2 Bd7
C19.21=Franskt:Winawer, 6...Ne7 7.Nf3 Nbc6 8.a4 Qa5+ 9.Bd2 Bd7 10.Bb5
C18.11=Franskt:Winawer, 6...Ne7 7.h4 Qc7 8.Nf3
C20.1=�ppet parti: 1.e4 e5
C20.2=�ppet parti: Mengarinis �ppning, 1.e4 e5 2.a3
C20.5=�ppet parti: 2.d3
C20.6=�ppet parti: 2.d3 d5
C20.3=�ppet parti: Patzer-Parnham �ppning, 1.e4 e5 2.Qh5
C20.4=�ppet parti: Napoleons �ppning, 1.e4 e5 2.Qf3
C20.7=�ppet parti: 2.c4
C20.8=�ppet parti: Lopez-Mcleod �ppning, 1.e4 e5 2.c3
C20.9=�ppet parti: Lopez-Mcleod, Lasa gambit, 1.e4 e5 2.c3 f5
C20.10=�ppet parti: Alapins �ppning, 1.e4 e5 2.Ne2
C20.11=�ppet parti: Alapins �ppning, 1.e4 e5 2.Ne2 Nf6
C20.12=�ppet parti: Portuguisisk �ppning, 1.e4 e5 2.Bb5
C20.13=�ppet parti: Portuguiskt 1.e4 e5 2.Bb5 Nf6
C20.14=�ppet parti: Portuguisisk gambit, 1.e4 e5 2.Bb5 Nf6 3.d4
C20.15=�ppet parti: Portuguisisk, 2...c6
C21.1=Centrumspel 1.e4 e5 2.d4
C21.2=Centrumspel Maroczys f�rsvar, 1.e4 e5 2.d4 d6
C21.3=Centrumspel Maroczys f�rsvar, 3.dxe5
C21.4=Centrumspel Maroczys f�rsvar, Philidors gambit, 1.e4 e5 2.d4 d6 3.dxe5 Bd7
C21.5=Centrumspel Dambytesvarianten, 1.e4 e5 2.d4 d6 3.dxe5 dxe5 4.Qxd8+
C21.6=Centrumspel 1.e4 e5 2.d4 exd4
C21.7=Centrumspel 3.Nf3
C21.8=Centrumspel Kieseritskyvarianten, 1.e4 e5 2.d4 exd4 3.Nf3 c5 4.Bc4 b5
C21.9=Centrumspel Halasz gambit, 1.e4 e5 2.d4 exd4 3.f4
C21.10=Dansk gambit: 1.e4 e5 2.d4 exd4 3.c3
C21.11=Dansk gambit: Svenonius f�rsvar, 1.e4 e5 2.d4 exd4 3.c3 Ne7
C21.12=Dansk gambit: S�rensens f�rsvar, 1.e4 e5 2.d4 exd4 3.c3 d5
C21.13=Dansk gambit: Antagen, 1.e4 e5 2.d4 exd4 3.c3 dxc3
C21.14=Dansk gambit: Antagen, 4.Bc4
C21.15=Dansk gambit: Antagen, 4.Bc4 cxb2 5.Bxb2
C21.16=Dansk gambit: K�penhamns f�rsvar, 2.d4 exd4 3.c3 dxc3 4.Bc4 cxb2 5.Bxb2 Bb4+
C21.17=Dansk gambit: Chigorins f�rsvar, 2.d4 exd4 3.c3 dxc3 4.Bc4 cxb2 5.Bxb2 Qe7
C21.18=Dansk gambit: Klassiskt f�rsvar, 2.d4 exd4 3.c3 dxc3 4.Bc4 cxb2 5.Bxb2 Nf6
C21.19=Dansk gambit: Schlechters f�rsvar, 2.d4 exd4 3.c3 dxc3 4.Bc4 cxb2 5.Bxb2 d5
C22.1=Centrumspel 1.e4 e5 2.d4 exd4 3.Qxd4
C22.2=Centrumspel 1.e4 e5 2.d4 exd4 3.Qxd4 Nc6
C22.3=Centrumspel Hallvarianten, 3.Qxd4 Nc6 4.Qc4
C22.4=Centrumspel Paulsen attack, 3.Qxd4 Nc6 4.Qe3
C22.5=Centrumspel Charousekvarianten, 3.Qxd4 Nc6 4.Qe3 Bb4+ 5.c3 Be7
C22.6=Centrumspel Bergervarianten, 3.Qxd4 Nc6 4.Qe3 Nf6
C22.7=Centrumspel Kupreichikvarianten, 3.Qxd4 Nc6 4.Qe3 Nf6 5.Nc3 Bb4 6.Bd2 O-O 7.O-O-O Re8 8.Bc4 d6 9.Nh3
C23.1=L�parspel 1.e4 e5 2.Bc4
C23.2=L�parspel Anderssens gambit
C23.3=L�parspel Philidors motattack
C23.4=L�parspel Lisitsins variant
C23.5=L�parspel Calabreses motgambit
C23.6=L�parspel Calabreses motgambit, J�nischvarianten
C23.7=L�parspel Klassiska varianten
C23.8=L�parspel 2...Bc5 3.Qe2
C23.9=L�parspel Lopez gambit
C23.10=L�parspel Lewis gambit
C23.11=L�parspel MacDonnells gambit
C23.12=L�parspel MacDonnells Dubbelgambit
C23.13=L�parspel MacDonnells, Fyra b�nder gambit
C23.14=L�parspel Philidorvarianten
C23.15=L�parspel del Rio-varianten
C23.16=L�parspel Lewis motgambit
C23.17=L�parspel Lewis motgambit, J�nisch
C23.18=L�parspel 2...Bc5 3.c3 Nf6
C23.19=L�parspel Prattvarianten
C24.1=L�parspel Berlin f�rsvar
C24.2=L�parspel Grecos gambit
C24.3=L�parspel 3.d3
C24.4=L�parspel 3.d3 d5
C24.5=L�parspel Paulsen f�rsvar
C24.6=L�parspel 3.d4
C24.7=L�parspel Urusovs gambit
C24.8=L�parspel Urusovs gambit, Panovvarianten
C24.9=L�parspel Urusovs gambit, Marshallvarianten
C24.10=L�parspel Urusovs gambit, 6.Bg5 Nc6 f�rsvar
C24.11=L�parspel Urusovs gambit, 7...c6 f�rsvar
C24.12=L�parspel Urusovs gambit, Larsenvarianten
C24.13=L�parspel Urusovs gambit, Karpovvarianten
C24.14=L�parspel Urusovs gambit, Forintos/Haagvarianten
C24.15=L�parspel Urusovs gambit, 7...Nc6 f�rsvar
C24.16=L�parspel Urusovs gambit, Keresvarianten
C24.17=L�parspel Urusovs gambit, Estrinvarianten
C25.1=Viennaparti
C25.2=Vienna: 2...Bb4
C25.3=Vienna: Zhuravlev
C25.4=Vienna: 2...d6
C25.5=Vienna: 2...d6 3.Bc4
C25.6=Vienna: 2...Bc5
C25.7=Vienna: Hammpe-Meitner
C25.8=Vienna: 2...Bc5 3.Bc4
C25.9=Vienna: 2...Bc5 3.Nf3
C25.10=Vienna: 2...Nc6
C25.11=Vienna: Fyfes gambit
C25.12=Vienna: Paulsenvarianten
C25.13=Vienna: Paulsen, 3...Bc5
C25.14=Vienna: 2...Nc6 3.Bc4
C25.15=Vienna: 2...Nc6 3.Bc4 Bc5
C25.16=Vienna: 2...Nc6 3.Bc4 Bc5 4.d3
C25.17=Vienna: 2...Nc6 3.Bc4 Bc5 4.Qg4
C25.18=Vienna: 2...Nc6 3.f4
C25.19=Vienna: 2...Nc6 3.f4
C25.20=Vienna: Steinitz gambit
C25.21=Vienna: Steinitz gambit, Fraser-Minckwitzvarianten
C25.22=Vienna: Steinitz gambit, Zukertort f�rsvar
C25.23=Vienna: 2...Nc6 3.f4 exf4 4.Nf3
C25.24=Vienna: 2...Nc6 3.f4 exf4 4.Nf3 g5
C25.25=Vienna: Hamppe-Muzios gambit
C25.26=Vienna: Hamppe-Muzio, Duboisvarianten
C25.27=Vienna: Hamppe-Allgaiers gambit
C25.28=Vienna: Hamppe-Allgaiers gambit, Alapinvarianten
C25.29=Vienna: Pierces gambit
C25.30=Vienna: Pierces gambit, Rushmere attack
C26.1=Vienna: 2...Nf6
C26.2=Vienna: Mengarinivarianten
C26.3=Vienna: 2...Nf6 3.d3
C26.4=Vienna: Smyslovvarianten
C26.5=Vienna: Smyslov, 3...Nc6
C26.6=Vienna: Smyslov, 3...Nc6
C26.7=Vienna: Smyslov, 3...Bc5
C26.8=Vienna: Smyslov, 3...Bc5
C26.9=Vienna: Smyslov, 3...Bc5 4.Bg2 d6
C26.10=Vienna: Smyslov, 3...Bc5 4.Bg2 O-O
C26.11=Vienna: Smyslov, 3...Bc5 4.Bg2 Nc6
C26.12=Vienna: Smyslov, 3...Bc5 4.Bg2 Nc6 5.Nge2
C26.13=Vienna: Smyslov, 3...d5
C26.14=Vienna: Smyslov, 3...d5
C26.15=Vienna: Smyslov, 3...d5, 5...Nxc3
C26.16=Vienna: Smyslov, 3...d5, 5...Nxc3 6.bxc3 Bd6
C26.17=Vienna: 3.Bc4
C26.18=Vienna: Horwitz gambit
C26.19=Vienna: 3.Bc4 Bb4
C26.20=Vienna: 3.Bc4 Bb4 4.Nf3
C26.21=Vienna: 3.Bc4 Bb4 4.Nf3 O-O
C26.22=Vienna: 3.Bc4 Bc5
C26.23=Vienna: 3.Bc4 Bc5 4.f4
C26.24=Vienna: 3.Bc4 Bc5 4.Nf3
C26.25=Vienna: 3.Bc4 Bc5 4.d3
C26.26=Vienna: 3.Bc4 Bc5 4.d3 d6
C26.27=Vienna: 3.Bc4 Bc5 4.d3 d6 5.Na4
C26.28=Vienna: 3.Bc4 Bc5 4.d3 d6 5.f4
C27.1=Vienna: 3.Bc4 Nxe4
C27.2=Vienna: 3.Bc4 Nxe4 4.Nxe4
C27.3=Vienna: 3.Bc4 Nxe4 4.Qh5
C27.4=Vienna: 3.Bc4 Nxe4 4.Qh5 Nd6 5.Qxe5+
C27.5=Vienna: 3.Bc4 Nxe4 4.Qh5 Nd6 5.Bb3
C27.6=Vienna: 3.Bc4 Nxe4 4.Qh5 Nd6 5.Bb3 Be7
C27.7=Vienna: Alekhinevarianten
C27.8=Vienna: 3.Bc4 Nxe4 4.Qh5 Nd6 5.Bb3 Nc6
C27.9=Vienna: Adams gambit
C27.10=Vienna: 3.Bc4 Nxe4 4.Qh5 Nd6 5.Bb3 Nc6
C27.11=Vienna: Frankenstein-Draculavarianten
C27.12=Vienna: Frankenstein-Dracula, 11.d3
C28.1=Vienna: 3.Bc4 Nc6
C28.2=Vienna: 3.Bc4 Nc6 4.f4
C28.3=Vienna: Bronsteins gambit
C28.4=Vienna: 3.Bc4 Nc6 4.d3
C28.5=Vienna: 3.Bc4 Nc6 4.d3 Be7
C28.6=Vienna: 3.Bc4 Nc6 4.d3 Na5
C28.7=Vienna: 3.Bc4 Nc6 4.d3 Na5 5.Nge2
C28.8=Vienna: 3.Bc4 Nc6 4.d3 Bc5
C28.9=Vienna: 3.Bc4 Nc6 4.d3 Bc5 5.Bg5
C28.10=Vienna: 3.Bc4 Nc6 4.d3 Bc5 5.f4
C28.11=Vienna: 3.Bc4 Nc6 4.d3 Bc5 5.f4 d6 6.Nf3
C28.12=Vienna: 3.Bc4 Nc6 4.d3 Bc5 5.f4 d6 6.Nf3 Bg4
C28.13=Vienna: 3.Bc4 Nc6 4.d3 Bc5 5.f4 d6 6.Nf3 a6
C28.14=Vienna: 3.Bc4 Nc6 4.d3 Bb4
C28.15=Vienna: 3.Bc4 Nc6 4.d3 Bb4 5.Nf3
C28.16=Vienna: 3.Bc4 Nc6 4.d3 Bb4 5.Bg5
C28.17=Vienna: 3.Bc4 Nc6 4.d3 Bb4 5.Ne2
C29.1=Vienna gambit
C29.2=Vienna gambit: 3...exf4
C29.3=Vienna gambit: 3...d6
C29.4=Vienna gambit: 3...d6 4.Nf3
C29.5=Vienna gambit: 3...d5
C29.6=Vienna gambit: 3...d5 4.exd5
C29.7=Vienna gambit: 3...d5 4.exd5 exf4
C29.8=Vienna gambit: Steinitzvarianten
C29.9=Vienna gambit: 4.fxe5
C29.10=Vienna gambit: 4.fxe5
C29.11=Vienna gambit: Oxfordvarianten
C29.12=Vienna gambit: Wurzburgers f�lla
C29.13=Vienna gambit: Oxford, 5...Bb4
C29.14=Vienna gambit: Oxford, 5...Bb4 6.dxe4 Qh4+ 7.Ke2
C29.15=Vienna gambit: Oxford, 5...Nxc3
C29.16=Vienna gambit: Oxford, 5...Nxc3 6.bxc3 d4
C29.17=Vienna gambit: Paulsen attack
C29.18=Vienna gambit: Paulsen attack, 5...Nc6
C29.19=Vienna gambit: Paulsen attack, Bardelebenvarianten
C29.20=Vienna gambit: Paulsen attack, Heydevarianten
C29.21=Vienna gambit: Paulsen attack, 5...Nxc3
C29.22=Vienna gambit: 5.Nf3
C29.23=Vienna gambit: 5.Nf3 Bg4
C29.24=Vienna gambit: Kaufmannvarianten
C29.25=Vienna gambit: 5.Nf3 Bb4
C29.26=Vienna gambit: 5.Nf3 Nc6
C29.27=Vienna gambit: Breyervarianten
C29.28=Vienna gambit: Breyer, 6.Qe2
C29.29=Vienna gambit: Breyer, 6.Qe2 Nxc3
C29.30=Vienna gambit: Breyer, 6.Qe2 Nxc3 7.dxc3
C30.1=Kungsgambit
C30.2=Kungsgambit: Mafias f�rsvar
C30.3=Kungsgambit: 2...d6
C30.4=Kungsgambit: 2...d6 3.Nf3
C30.5=Kungsgambit: 2...d6 3.Nf3 Nc6
C30.6=Kungsgambit: Wadevarianten
C30.7=Kungsgambit: Norwaldvarianten
C30.8=Kungsgambit: Norwaldvarianten, Schubert line
C30.9=Kungsgambit: Norwaldvarianten, B�cker gambit
C30.10=Kungsgambit: Keene f�rsvar
C30.11=Kungsgambit: Keene f�rsvar, 3.g3 Qe7
C30.12=Kungsgambit: 2...Nc6
C30.13=Kungsgambit: Adelaide-Wahlsvarianten
C30.14=Kungsgambit: Adelaide-Wahls, 4.exf5
C30.15=Kungsgambit: Adelaide-Wahls, 4.exf5 e4
C30.16=Kungsgambit: Adelaide-Wahls, 4.exf5 e4 5.Ne5 Nf6
C30.17=Kungsgambit: Avb�jd Klassisk kungsgambit
C30.18=Avb�jd Kungsgambit Klassisk, 3.Bc4
C30.19=Avb�jd Kungsgambit Klassisk, 3.Nf3
C30.20=Avb�jd Kungsgambit Klassisk, Senechauds motgambit
C30.21=Avb�jd Kungsgambit Klassisk, 3.Nf3 d6
C30.22=Avb�jd Kungsgambit Klassisk, Heathvarianten
C30.23=Avb�jd Kungsgambit Klassisk, Soldatenkov-varianten
C30.24=Avb�jd Kungsgambit Klassisk, 3.Nf3 d6 4.Nc3
C30.25=Avb�jd Kungsgambit Klassisk, Hanhamvarianten
C30.26=Avb�jd Kungsgambit Klassisk, 3.Nf3 d6 4.Nc3 Nf6 5.Bc4
C30.27=Avb�jd Kungsgambit Klassisk, Svenonius-varianten
C30.28=Avb�jd Kungsgambit Klassisk, 4.c3
C30.29=Avb�jd Kungsgambit Klassisk, Marshall attack
C30.30=Avb�jd Kungsgambit Klassisk, 4.c3 Bb6
C30.31=Avb�jd Kungsgambit Klassisk, 4.c3 Nf6
C30.32=Avb�jd Kungsgambit Klassisk, 4.c3 Nf6 5.d4
C30.33=Avb�jd Kungsgambit Klassisk, 4.c3 Nf6 5.d4
C30.34=Avb�jd Kungsgambit Klassisk, 4.c3 Nf6 5.d4
C30.35=Avb�jd Kungsgambit Klassisk motgambit
C30.36=Avb�jd Kungsgambit Klassisk, Retisvarianten
C31.1=Avb�jd Kungsgambit Falkbeers motgambit
C31.2=Avb�jd Kungsgambit Falkbeer, Tartakowervarianten
C31.3=Avb�jd Kungsgambit Falkbeer, Milner-Barryvarianten
C31.4=Avb�jd Kungsgambit Falkbeer, 3.exd5
C31.5=Avb�jd Kungsgambit Falkbeer, 3.exd5 exf4
C31.6=Avb�jd Kungsgambit Falkbeer, Marshall/Nimzowitsch motgambit
C31.7=Avb�jd Kungsgambit Falkbeer, Marshall/Nimzowitsch, 4.dxc6
C31.8=Avb�jd Kungsgambit Falkbeer, Marshall/Nimzowitsch, 4.Qe2
C31.9=Avb�jd Kungsgambit Falkbeer, Marshall/Nimzowitsch, 4.Nc3
C31.10=Avb�jd Kungsgambit Falkbeer, 3.exd5 e4
C31.11=Avb�jd Kungsgambit Falkbeer, Rubinsteinvarianten
C31.12=Avb�jd Kungsgambit Falkbeer, Nimzowitschvarianten
C31.13=Avb�jd Kungsgambit Falkbeer, 4.d3
C32.1=Avb�jd Kungsgambit Falkbeer, 4.d3 Nf6
C32.2=Avb�jd Kungsgambit Falkbeer, Keresvarianten
C32.3=Avb�jd Kungsgambit Falkbeer, Keres, 5...exd3
C32.4=Avb�jd Kungsgambit Falkbeer, Retisvarianten
C32.5=Avb�jd Kungsgambit Falkbeer, 4.d3 Nf6 5.Nc3
C32.6=Avb�jd Kungsgambit Falkbeer, 4.d3 Nf6 5.Nc3 Bb4
C32.7=Avb�jd Kungsgambit Falkbeer, Morphy gambit
C32.8=Avb�jd Kungsgambit Falkbeer, 5.dxe4
C32.9=Avb�jd Kungsgambit Falkbeer, Charousekvarianten
C32.10=Avb�jd Kungsgambit Falkbeer, 5.dxe4 Nxe4 6.Be3
C32.11=Avb�jd Kungsgambit Falkbeer, 5.dxe4 Nxe4 6.Nf3
C32.12=Avb�jd Kungsgambit Falkbeer, 5.dxe4 Nxe4 6.Nf3 Bc5 7.Qe2
C32.13=Avb�jd Kungsgambit Falkbeer, Alapinvarianten
C32.14=Avb�jd Kungsgambit Falkbeer, Huvudvarianten, 7...Bf5
C32.15=Avb�jd Kungsgambit Falkbeer, Tarraschvarianten
C32.16=Avb�jd Kungsgambit Falkbeer, Huvudvarianten, 7...Bf5 8.Nc3
C33.1=Antagen Kungsgambit
C33.2=Antagen Kungsgambit: Tumbleweed/Drunken King
C33.3=Antagen Kungsgambit: Orsinis gambit
C33.4=Antagen Kungsgambit: Stammas (Leonardo) gambit
C33.5=Antagen Kungsgambit: Schurigs gambit
C33.6=Antagen Kungsgambit: Basmans gambit
C33.7=Antagen Kungsgambit: Carreras gambit
C33.8=Antagen Kungsgambit: Eisenbergs gambit
C33.9=Antagen Kungsgambit: Eisenbergs gambit
C33.10=Antagen Kungsgambit: Villemsons gambit
C33.11=Antagen Kungsgambit: Keres gambit
C33.12=Antagen Kungsgambit: Breyers gambit
C33.13=Antagen Kungsgambit: Mindre l�pares (Tartakower) gambit
C33.14=Antagen Kungsgambit: L�pargambit
C33.15=Antagen Kungsgambit: L�pargambit, Chigorins attack
C33.16=Antagen Kungsgambit: L�pargambit, Grecovarianten
C33.17=Antagen Kungsgambit: L�pargambit, Klassiskt f�rsvar
C33.18=Antagen Kungsgambit: L�pargambit, Grimms attack
C33.19=Antagen Kungsgambit: L�pargambit, Klassiskt f�rsvar
C33.20=Antagen Kungsgambit: L�pargambit, McDonnells attack
C33.21=Antagen Kungsgambit: bishop's gambit, McDonnells attack
C33.22=Antagen Kungsgambit: L�pargambit, Fraservarianten
C33.23=Antagen Kungsgambit: L�pargambit, Klassisk f�rsvar, Cozio attack
C33.24=Antagen Kungsgambit: L�pargambit, Bodens f�rsvar
C33.25=Antagen Kungsgambit: L�pargambit, Bryans motgambit
C33.26=Antagen Kungsgambit: L�pargambit, Bryans motgambit
C33.27=Antagen Kungsgambit: L�pargambit, Steinitz f�rsvar
C33.28=Antagen Kungsgambit: L�pargambit, Maurian f�rsvar
C33.29=Antagen Kungsgambit: L�pargambit, Ruy Lopez f�rsvar
C33.30=Antagen Kungsgambit: L�pargambit, Lopez-Gianutios motgambit
C33.31=Antagen Kungsgambit: L�pargambit, Lopez-Gianutios motgambit, Heinvarianten
C33.32=Antagen Kungsgambit: L�pargambit, Bledowvarianten
C33.33=Antagen Kungsgambit: L�pargambit, Bledow, 4.exd5
C33.34=Antagen Kungsgambit: L�pargambit, Bledow, 4.Bxd5
C33.35=Antagen Kungsgambit: L�pargambit, Boren-Svenoniusvarianten
C33.36=Antagen Kungsgambit: L�pargambit, Anderssenvarianten
C33.37=Antagen Kungsgambit: L�pargambit, Morphyvarianten
C33.38=Antagen Kungsgambit: L�pargambit, Cozio f�rsvar
C33.39=Antagen Kungsgambit: L�pargambit, Bogoljubowvarianten
C33.40=Antagen Kungsgambit: L�pargambit, Paulsens attack
C33.41=Antagen Kungsgambit: L�pargambit, J�nischvarianten
C34.1=Antagen Kungsgambit: King's Knight gambit
C34.2=Antagen Kungsgambit: Bonsch-Osmolovskyvarianten
C34.3=Antagen Kungsgambit: Gianutios motgambit
C34.4=Antagen Kungsgambit: Beckers f�rsvar (Anti-Kieseritzky)
C34.5=Antagen Kungsgambit: Schallops f�rsvar
C34.6=Antagen Kungsgambit: Fischers f�rsvar
C34.7=Antagen Kungsgambit: Fischer, 4.Bc4
C34.8=Antagen Kungsgambit: Fischer, 4.d4
C34.9=Antagen Kungsgambit: Fischer, Huvudvarianten
C35.1=Antagen Kungsgambit: Cunninghams f�rsvar
C35.2=Antagen Kungsgambit: Cunningham, Bertins gambit
C35.3=Antagen Kungsgambit: Cunningham, Trebondegambit
C35.4=Antagen Kungsgambit: Cunningham, Euwes f�rsvar
C36.1=Antagen Kungsgambit: Skandinavisk (Abbazia)varianten
C36.2=Antagen Kungsgambit: Skandinavisk, 4.exd5
C36.3=Antagen Kungsgambit: Skandinavisk, 4.exd5 Bd6
C36.4=Antagen Kungsgambit: Skandinavisk, Moderna Varianten
C36.5=Antagen Kungsgambit: Skandinavisk, Modern, 5.Bc4
C36.6=Antagen Kungsgambit: Skandinavisk, Modern, 5.Nc3
C36.7=Antagen Kungsgambit: Skandinavisk, Modern, 5.Bb5+ 
C36.8=Antagen Kungsgambit: Skandinavisk, Modern, 5.Bb5+ c6
C36.9=Antagen Kungsgambit: Skandinavisk, Modern, 5.Bb5+ c6 6.dxc6 Nxc6
C36.10=Antagen Kungsgambit: Skandinavisk, Modern, 5.Bb5+ c6 6.dxc6 bxc6
C36.11=Antagen Kungsgambit: Skandinavisk, Botvinnikvarianten
C37.1=Antagen Kungsgambit: 3.Nf3 g5
C37.2=Antagen Kungsgambit: Quaades gambit
C37.3=Antagen Kungsgambit: Rosentreters gambit
C37.4=Antagen Kungsgambit: S�rensens gambit
C37.5=Antagen Kungsgambit: 3.Nf3 g5 4.Bc4
C37.6=Antagen Kungsgambit: Blachlys gambit
C37.7=Antagen Kungsgambit: 3.Nf3 g5 4.Bc4 g4
C37.8=Antagen Kungsgambit: Lollis gambit (Vild Muzio)
C37.9=Antagen Kungsgambit: Lollis gambit, Young-varianten
C37.10=Antagen Kungsgambit: Ghulam-Kassims gambit
C37.11=Antagen Kungsgambit: MacDonnells gambit
C37.12=Antagen Kungsgambit: Salvios gambit
C37.13=Antagen Kungsgambit: Salvio, Silberschmidts gambit
C37.14=Antagen Kungsgambit: Salvio, Anderssens motattack
C37.15=Antagen Kungsgambit: Salvio, Cochranes gambit
C37.16=Antagen Kungsgambit: Salvio, Herzfelds gambit
C37.17=Antagen Kungsgambit: Muzios gambit
C37.18=Antagen Kungsgambit: Muzios gambit, Paulsenvarianten
C37.19=Antagen Kungsgambit: Dubbel Muzios gambit
C37.20=Antagen Kungsgambit: Muzios gambit, Froms f�rsvar
C37.21=Antagen Kungsgambit: Muzios gambit, Holloways f�rsvar
C37.22=Antagen Kungsgambit: Muzios gambit, Kling and Horwitz motattack
C37.23=Antagen Kungsgambit: Muzios gambit, Brentanos f�rsvar
C38.1=Antagen Kungsgambit: 3.Nf3 g5 4.Bc4 Bg7
C38.2=Antagen Kungsgambit: Hansteins gambit
C38.3=Antagen Kungsgambit: Hansteins gambit
C38.4=Antagen Kungsgambit: Philidors gambit
C38.5=Antagen Kungsgambit: Grecos gambit
C38.6=Antagen Kungsgambit: Philidors gambit, Schultzvarianten
C39.1=Antagen Kungsgambit: 3.Nf3 g5 4.h4
C39.2=Antagen Kungsgambit: Allgaiers gambit
C39.3=Antagen Kungsgambit: Allgaiers,Hornys f�rsvar
C39.4=Antagen Kungsgambit: Allgaier, Thoroldvarianten
C39.5=Antagen Kungsgambit: Allgaier, Cookvarianten
C39.6=Antagen Kungsgambit: Allgaier, Blackburnes gambit
C39.7=Antagen Kungsgambit: Allgaier, Walkers attack
C39.8=Antagen Kungsgambit: Allgaier, Urusovs attack
C39.9=Antagen Kungsgambit: Allgaier, Schlechters f�rsvar
C39.10=Antagen Kungsgambit: Kieseritsky
C39.11=Antagen Kungsgambit: Kieseritsky, Greenvarianten
C39.12=Antagen Kungsgambit: Kieseritsky, Paulsen f�rsvar
C39.13=Antagen Kungsgambit: Kieseritsky, Long Whip f�rsvar
C39.14=Antagen Kungsgambit: Kieseritsky, Long Whip f�rsvar, J�nischvarianten
C39.15=Antagen Kungsgambit: Kieseritsky, Brentanos (Campbell) f�rsvar
C39.16=Antagen Kungsgambit: Kieseritsky, Brentanos f�rsvar, Kaplanekvarianten
C39.17=Antagen Kungsgambit: Kieseritsky, Brentanos f�rsvar
C39.18=Antagen Kungsgambit: Kieseritsky, Brentanos f�rsvar, Carovarianten
C39.19=Antagen Kungsgambit: Kieseritsky, Salvios (Rosenthal) f�rsvar
C39.20=Antagen Kungsgambit: Kieseritsky, Salvios f�rsvar, Coziovarianten
C39.21=Antagen Kungsgambit: Kieseritsky, Polerios f�rsvar
C39.22=Antagen Kungsgambit: Kieseritsky, Neumanns f�rsvar
C39.23=Antagen Kungsgambit: Kieseritsky, Berlinf�rsvaret
C39.24=Antagen Kungsgambit: Kieseritsky, Berlinf�rsvaret, Rivierevarianten
C39.25=Antagen Kungsgambit: Kieseritsky, Berlinf�rsvaret, 6.Bc4
C39.26=Antagen Kungsgambit: Kieseritsky, Rice gambit
C40.1=�ppet parti
C40.2=�ppet parti: Damianos f�rsvar
C40.3=�ppet parti: Grecos f�rsvar
C40.4=�ppet parti: Gunderams f�rsvar
C40.5=Elefantgambit
C40.6=Elefantgambit: 3.Nxe5
C40.7=Elefantgambit: 3.Nxe5 dxe4 4.Bc4
C40.8=Elefantgambit: 3.exd5
C40.9=Elefantgambit: Maroczy
C40.10=Elefantgambit: Paulsen
C40.11=Lettisk gambit
C40.12=Lettisk gambit: 3.d3
C40.13=Lettisk gambit: 3.Nc3
C40.14=Lettisk gambit: 3.d4
C40.15=Lettisk gambit: 3.d4 fxe4 5.Nxe5 Nf6
C40.16=Lettisk gambit: 3.exf5
C40.17=Lettisk gambit: 3.exf5 e4
C40.18=Lettisk gambit: 3.Bc4
C40.19=Lettisk gambit: Strautinsvarianten
C40.20=Lettisk gambit: Morgadovarianten
C40.21=Lettisk gambit: 3.Bc4 fxe4
C40.22=Lettisk: Blackburnevarianten (Corkscrew motgambit)
C40.23=Lettisk gambit: Svedenborgvarianten
C40.24=Lettisk gambit: Svedenborg, 6.Nxg6 Nf6
C40.25=Lettisk gambit: Svedenborg, 6.Nxg6 hxg6
C40.26=Lettisk gambit: F�rgiftad bonde-varianten
C40.27=Lettisk gambit: F�rgiftad bonde, Huvudvarianten
C40.28=Lettisk gambit: 3.Nxe5
C40.29=Lettisk gambit: 3.Nxe5 Nc6
C40.30=Lettisk gambit: 3.Nxe5 Qf6
C40.31=Lettisk gambit: 3.Nxe5 Qf6 4.Nc4
C40.32=Lettisk gambit: 3.Nxe5 Qf6 4.d4
C40.33=Lettisk gambit: 3.Nxe5 Qf6 4.d4 d6
C40.34=Lettisk gambit: 3.Nxe5 Qf6 4.d4 d6 5.Nc4
C40.35=Lettisk gambit: 3.Nxe5 Qf6 4.d4 d6 5.Nc4 fxe4
C40.36=Lettisk gambit: 3.Nxe5 Qf6 4.d4 d6 5.Nc4 fxe4 6.Be2
C40.37=Lettisk gambit: Nimzowitschvarianten
C40.38=Lettisk gambit: 3.Nxe5 Qf6 4.d4 d6 5.Nc4 fxe4 6.Nc3
C41.1=Philidors f�rsvar
C41.2=Philidor: 3.Bc4
C41.3=Philidor: Steinitzvarianten
C41.4=Philidor: Lopez motgambit
C41.5=Philidor: Lopez motgambit, J�nischvarianten
C41.6=Philidor: 3.d4
C41.7=Philidor: Philidors motgambit
C41.8=Philidor: Philidors motgambit, Zukertortvarianten
C41.9=Philidor: Philidors motgambit, 4.dxe5
C41.10=Philidor: Philidors motgambit, Steinitzvarianten
C41.11=Philidor: Philidors motgambit, del Rio attack
C41.12=Philidor: Philidors motgambit, Bergervarianten
C41.13=Philidor: Hanhamvarianten
C41.14=Philidor: Hanham, 4.Bc4
C41.15=Philidor: Hanham, 4.Bc4 c6
C41.16=Philidor: Hanham, Krausevarianten
C41.17=Philidor: Hanham, Steinervarianten
C41.18=Philidor: Hanham, Kmochvarianten
C41.19=Philidor: Hanham, Bergervarianten
C41.20=Philidor: Hanham, Schlechtervarianten
C41.21=Philidor: Hanham, Delmarvarianten
C41.22=Philidor: 3...exd4
C41.23=Philidor: Birds gambit
C41.24=Philidor: Morphyvarianten
C41.25=Philidor: Morphy, 4...Nc6
C41.26=Philidor: Morphy, 4...Nf6
C41.27=Philidor: Morphy, 4...Nf6 5.Nc3
C41.28=Philidor: 3...exd4 4.Nxd4
C41.29=Philidor: Paulsen attack
C41.30=Philidor: 3...exd4 4.Nxd4 Nf6
C41.31=Philidor: 3...exd4 4.Nxd4 Nf6 5.Nc3
C41.32=Philidor: 3...exd4 4.Nxd4 Nf6 5.Nc3 Be7
C41.33=Philidor: 3...exd4 4.Nxd4 Nf6 5.Nc3 Be7 6.Bc4
C41.34=Philidor: Antoshinvarianten
C41.35=Philidor: Bergervarianten
C41.36=Philidor: Larsenvarianten
C41.37=Philidor: Nimzowitschvarianten
C41.38=Philidor: Nimzowitsch, Kleinvarianten
C41.39=Philidor: Nimzowitsch, Locockvarianten
C41.40=Philidor: Avbytesvarianten
C41.41=Philidor: Avbyte, Sokolskyvarianten
C41.42=Philidor: Avbyte, Rellstabvarianten
C41.43=Philidor: Nimzowitschvarianten
C41.44=Philidor: F�rb�ttrad Hanham
C41.45=Philidor: F�rb�ttrad Hanham, 5.Bc4
C41.46=Philidor: F�rb�ttrad Hanham, 5.Bc4 Be7
C41.47=Philidor: F�rb�ttrad Hanham, 6.Bxf7+
C41.48=Philidor: F�rb�ttrad Hanham, 6.Ng5
C41.49=Philidor: F�rb�ttrad Hanham, Larobokvarianten
C41.50=Philidor: F�rb�ttrad Hanham, 6.dxe5
C41.51=Philidor: F�rb�ttrad Hanham, 6.dxe5 Nxe5
C41.52=Philidor: F�rb�ttrad Hanham, 6.dxe5 dxe5
C41.53=Philidor: F�rb�ttrad Hanham 6.O-O
C41.54=Philidor: F�rb�ttrad Hanham, Huvudvarianten
C41.55=Philidor: F�rb�ttrad Hanham, 7.a4
C41.56=Philidor: F�rb�ttrad Hanham, 7.a4 c6
C41.57=Philidor: F�rb�ttrad Hanham, 7.Qe2
C41.58=Philidor: F�rb�ttrad Hanham, 7.Qe2 c6 8.a4
C41.59=Philidor: F�rb�ttrad Hanham, Sozinvarianten
C41.60=Philidor: F�rb�ttrad Hanham, 7.Re1
C41.61=Philidor: F�rb�ttrad Hanham, 7.Re1 c6 8.a4
C41.62=Philidor: F�rb�ttrad Hanham, 7.Re1 c6 8.a4 b6
C42.1=Ryskt parti (Petroffs f�rsvar)
C42.2=Ryskt parti: 3.d3
C42.3=Ryskt-Trespringar parti
C42.4=Ryskt-Trespringar parti
C42.5=Ryskt-Trespringar parti, 4.Nxe5
C42.6=Ryskt parti: Italiensk variant
C42.7=Ryskt parti: Boden-Kieseritskys gambit
C42.8=Ryskt parti: Antagen Boden-Kieseritskys gambit
C42.9=Ryskt parti: 3.Nxe5
C42.10=Ryskt parti: Damianovarianten
C42.11=Ryskt parti: 3.Nxe5 d6
C42.12=Ryskt parti: Cochranes gambit
C42.13=Ryskt parti: Cochranes gambit, 5.d4
C42.14=Ryskt parti: Paulsens attack
C42.15=Ryskt parti: 3.Nxe5 d6 4.Nf3
C42.16=Ryskt parti: Fransk attack
C42.17=Ryskt parti: Vienna/Kaufmann
C42.18=Ryskt parti: Nimzowitsch attack
C42.19=Ryskt parti: Cozio/Lasker
C42.20=Ryskt parti: Milner-Barryvarianten
C42.21=Ryskt parti: 5.Qe2, Dambyte
C42.22=Ryskt parti: Klassisk
C42.23=Ryskt parti: Klassisk, St�ngd variant
C42.24=Ryskt parti: Klassisk, 5...d5
C42.25=Ryskt parti: Klassisk, 6.Bd3
C42.26=Ryskt parti: Klassisk, Marshallvarianten
C42.27=Ryskt parti: Klassisk, Tarraschvarianten
C42.28=Ryskt parti: Klassisk, Marshalls f�lla
C42.29=Ryskt parti: Klassisk, Marshall, 8.c4 c6
C42.30=Ryskt parti: Klassisk, 6.Bd3 Be7
C42.31=Ryskt parti: Klassisk, Masonvarianten
C42.32=Ryskt parti: Klassisk, 6.Bd3 Be7 7.O-O Nc6
C42.33=Ryskt parti: Klassisk, J�nischvarianten
C42.34=Ryskt parti: Klassisk, J�nisch, Huvudvarianten
C42.35=Ryskt parti: Klassisk, Chigorinvarianten
C42.36=Ryskt parti: Klassisk, Chigorin, 8...Bf5
C42.37=Ryskt parti: Klassisk, Chigorin, 8...Bg4
C42.38=Ryskt parti: Klassisk, Chigorin, 8...Bg4 9.c4
C42.39=Ryskt parti: Klassisk, Chigorin, 8...Bg4 9.c3
C42.40=Ryskt parti: Klassisk, Bergervarianten
C42.41=Ryskt parti: Klassisk, Krausevarianten
C42.42=Ryskt parti: Klassisk, Maroczyvarianten
C43.1=Ryskt parti: Moderna (Steinitz) attack
C43.2=Ryskt parti: Modern attack
C43.3=Ryskt parti: Modern attack
C43.4=Ryskt parti: Modern attack, Tals gambit
C43.5=Ryskt parti: Modern attack, Steinitzvarianten
C43.6=Ryskt parti: Modern attack, Bardelebenvarianten
C43.7=Ryskt parti: Modern attack, 3...exd4, Huvudvarianten
C43.8=Ryskt parti: Modern attack, 3...exd4, Huvudvarianten, 7.Nc3
C43.9=Ryskt parti: Modern attack, Pillsburyvarianten
C43.10=Ryskt parti: Modern attack, 3...Nxe4
C43.11=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3
C43.12=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 Nc6
C43.13=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 Nc6 5.d5
C43.14=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 Nc6 5.Bxe4
C43.15=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5
C43.16=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.dxe5
C43.17=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5
C43.18=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5 Nc6
C43.19=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5 Be7
C43.20=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5 Bd6
C43.21=Ryskt parti: Modern attack, Trifunovicvarianten
C43.22=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5 Nd7
C43.23=Ryskt parti: Modern attack, 3...Nxe4 4.Bd3 d5 5.Nxe5 Nd7 6.Nxd7
C43.24=Ryskt parti: Modern attack, 3...Nxe4, Huvudvarianten
C43.25=Ryskt parti: Modern attack, 3...Nxe4, Huvudvarianten, 7...Qh4
C43.26=Ryskt parti: Modern attack, 3...Nxe4, Huvudvarianten, 7...Bd6
C44.1=�ppet parti
C44.2=�ppet parti: Irl�ndsk (Chicago) gambit
C44.3=�ppet parti: Paschmans vingambit
C44.4=�ppet parti: Dresden�ppning
C44.5=�ppet parti: Konstantinopolsky
C44.6=�ppet parti: Inverterad Ungersk
C44.7=�ppet parti: Taylers �ppning
C44.8=�ppet parti: Inverterad Philidor
C44.9=�ppet parti: Inverterad Philidor
C44.10=�ppet parti: Inverterad Philidor
C44.11=�ppet parti: Inverterad Philidor, 4.g3
C44.12=�ppet parti: Inverterad Philidor, 4.Be2
C44.13=�ppet parti: Inverterad Hanham
C44.14=Ponzianis �ppning
C44.15=Ponziani: Retisvarianten
C44.16=Ponziani: Romanishinvarianten
C44.17=Ponzianis motgambit
C44.18=Ponzianis motgambit, Schmidtattacken
C44.19=Ponzianis motgambit, Cordelvarianten
C44.20=Ponziani: 3...d5
C44.21=Ponziani: 3...d5 4.Qa4
C44.22=Ponziani: Carovarianten
C44.23=Ponziani: Leonhardtvarianten
C44.24=Ponziani: Steinitzvarianten
C44.25=Ponziani: 3...Nf6
C44.26=Ponziani: 3...Nf6
C44.27=Ponziani: 3...Nf6 4.d4 exd4
C44.28=Ponziani: 3...Nf6 4.d4 Nxe4
C44.29=Ponziani: Frasers f�rsvar
C44.30=Ponziani: 3...Nf6 4.d4 Nxe4 5.d5 Ne7
C44.31=Skottsk �ppning
C44.32=Skottskt: Lollivarianten
C44.33=Skottskt: Cochranevarianten
C44.34=Skottskt: 3...d6
C44.35=Skottskt: 3...exd4
C44.36=Skottskt: Relfssons gambit
C44.37=Skottskt: G�ringgambit
C44.38=Skottskt: G�ringgambit, 4...d5
C44.39=Skottskt: G�ringgambit, 4...d3
C44.40=Skottskt: G�ringgambit, 4...dxc3
C44.41=Skottskt: G�ringgambit, 4...dxc3 5.Bc4
C44.42=Skottskt: G�ringgambit, 4...dxc3 5.Bc4 cxb2 6.Bxb2
C44.43=Skottskt: G�ringgambit, 4...dxc3 5.Nxc3
C44.44=Skottskt: G�ringgambit, 4...dxc3 5.Nxc3 Bb4
C44.45=Skottskt: G�ringgambit, Bardelebenvarianten
C44.46=Skottskt: G�ringgambit, 4...dxc3 5.Nxc3 Bb4 6.Bc4 d6
C44.47=Skottskt: G�ringgambit, 4...dxc3 5.Nxc3 Bb4 6.Bc4 d6 7.O-O
C44.48=Skottsk gambit
C44.49=Skottsk gambit: London f�rsvar
C44.50=Skottsk gambit: 4...Bc5
C44.51=Skottsk gambit: 5.Ng5
C44.52=Skottsk gambit: Vitzhums attack
C44.53=Skottsk gambit: 5.O-O
C44.54=Skottsk gambit: Anderssens (Paulsen) motattack
C44.55=Skottsk gambit: 5.c3
C44.56=Skottsk gambit: 5.c3 d3
C45.1=Skottskt: 4.Nxd4
C45.2=Skottskt: 4.Nxd4 Nxd4
C45.3=Skottskt: Ghulam Kassimvarianten
C45.4=Skottskt: 4.Nxd4 Bb4+
C45.5=Skottskt: 4.Nxd4 Qf6
C45.6=Skottskt: Steinitzvarianten
C45.7=Skottskt: Steinitz, 5.Qd3
C45.8=Skottskt: Steinitz, Fraser attack
C45.9=Skottskt: Steinitz, 5.Nc3
C45.10=Skottskt: Steinitz, 5.Nb5
C45.11=Skottskt: Steinitz, 5.Nb5 Qxe4+
C45.12=Skottskt: Steinitz, 5.Nb5 Bc5
C45.13=Skottskt: Steinitz, 5.Nb5 Bc5 6.Qf3
C45.14=Skottskt: Steinitz, 5.Nb5 Bb4+
C45.15=Skottskt: Steinitz, Bergervarianten
C45.16=Skottskt: Steinitz, 5.Nb5 Bb4+ 6.Bd2
C45.17=Skottskt: Steinitz, Rosenthalvarianten
C45.18=Skottskt: 4.Nxd4 Nf6
C45.19=Skottskt: 4.Nxd4 Nf6 5.Nxc6
C45.20=Skottskt: Tartakowervarianten
C45.21=Skottskt: 4.Nxd4 Nf6 5.Nxc6 bxc6 6.Bd3
C45.22=Skottskt: Miesesvarianten
C45.23=Skottskt: Mieses, 6...Qe7
C45.24=Skottskt: Mieses, 6...Qe7 7.Qe2
C45.25=Skottskt: Mieses, 8.c4
C45.26=Skottskt: Mieses, 8.c4 Ba6
C45.27=Skottskt: Mieses, 8.c4 Ba6 9.b3
C45.28=Skottskt: 4.Nxd4 Bc5
C45.29=Skottskt: 4.Nxd4 Bc5 5.Nb3
C45.30=Skottskt: Romanishinvarianten
C45.31=Skottskt: 4.Nxd4 Bc5 5.Nb3 Bb6
C45.32=Skottskt: 4.Nxd4 Bc5 5.Nb3 Bb6 6.a4
C45.33=Skottskt: 4.Nxd4 Bc5 5.Nb3 Bb6 6.a4 a6
C45.34=Skottskt: 4.Nxd4 Bc5 5.Nb3 Bb6 6.a4 a6 7.Nc3
C45.35=Skottskt: Gellervarianten
C45.36=Skottskt: 4.Nxd4 Bc5 5.Nb3 Bb6 6.a4 a6 7.Nc3 Qf6
C45.37=Skottskt: 4.Nxd4 Bc5 5.Nxc6
C45.38=Skottskt: 4.Nxd4 Bc5 5.Nxc6 Qf6 6.Qd2
C45.39=Skottskt: 4.Nxd4 Bc5 5.Nxc6 Qf6 6.Qd2 dxc6 7.Nc3
C45.40=Skottskt: 4.Nxd4 Bc5 5.Be3
C45.41=Skottskt: Blumenfeld attack
C45.42=Skottskt: 4.Nxd4 Bc5 5.Be3 Qf6 6.c3
C45.43=Skottskt: 4.Nxd4 Bc5 5.Be3 Qf6 6.c3 Nge7
C45.44=Skottskt: Blackburnes attack
C45.45=Skottskt: Meitnervarianten
C45.46=Skottskt: Paulsens attack
C45.47=Skottskt: Paulsen, Gunsbergs f�rsvar
C45.48=Skottskt: 4.Nxd4 Bc5 5.Be3 Qf6 6.c3 Nge7 7.Bc4
C45.49=Skottskt: 4.Nxd4 Bc5 5.Be3 Qf6 6.c3 Nge7 7.Bc4 Ne5
C46.1=Trespringar parti
C46.2=Trespringar: Winawers f�rsvar
C46.3=Trespringar: 3...d6
C46.4=Trespringar: 3...d6 4.d4
C46.5=Trespringar: 3...Bc5
C46.6=Trespringar: 3...Bc5 4.Bb5
C46.7=Trespringar: 3...Bc5 4.Nxe5
C46.8=Trespringar: 3...Bb4
C46.9=Trespringar: 3...Bb4 4.Nd5
C46.10=Trespringar: Schlechtervarianten
C46.11=Trespringar: Steinitzvarianten
C46.12=Trespringar: Steinitz, 4.d4
C46.13=Trespringar: Steinitz, Rosenthalvarianten
C46.14=Trespringar: Steinitz, 4.d4 exd4 5.Nxd4
C46.15=Trespringar: Steinitz, 4.d4 exd4 5.Nxd4 Bg7
C46.16=Trespringar: Steinitz, 4.d4 exd4 5.Nxd4 Bg7 6.Be3
C46.17=Trespringar: Steinitz, 4.d4 exd4 5.Nxd4 Bg7 6.Be3 Nf6
C47.1=Fyrspringarparti
C47.2=Fyra Springare: Halloween gambit
C47.3=Fyra Springare: Gunsbergvarianten
C47.4=Fyra Springare: Van der Wiel-varianten
C47.5=Fyra Springare: Italiensk variant
C47.6=Fyra Springare: Glekvarianten
C47.7=Fyra Springare: Glek, 4...d5
C47.8=Fyra Springare: Glek, 4...Bc5
C47.9=Fyra Springare: Glek, 4...Bc5
C47.10=Fyra Springare: Glek, Huvudvarianten
C47.11=Fyra Springare: Skottska Varianten
C47.12=Fyra Springare: Skottsk, 4...d6
C47.13=Fyra Springare: Skottsk, Bogoljubow
C47.14=Fyra Springare: Skottsk, Bogoljubow, 5.d5
C47.15=Fyra Springare: Skottsk, Krausevarianten
C47.16=Fyra Springare: Skottsk, 4...exd4
C47.17=Fyra Springare: Belgradgambit
C47.18=Fyra Springare: Belgradgambit, 5...Nb4
C47.19=Fyra Springare: Belgradgambit, 5...Nxd5
C47.20=Fyra Springare: Belgradgambit, 5...Nxe4
C47.21=Fyra Springare: Belgradgambit, 5...Nxe4 6.Qe2 (Gamla Line)
C47.22=Fyra Springare: Belgradgambit, 5...Nxe4 6.Bc4 (Moderna Line)
C47.23=Fyra Springare: Belgradgambit, 5...Be7
C47.24=Fyra Springare: Skottsk, 4...exd4 5.Nxd4
C47.25=Fyra Springare: Skottsk, 4...exd4 5.Nxd4 d6
C47.26=Fyra Springare: Skottsk, 4...exd4 5.Nxd4 Bc5
C47.27=Fyra Springare: Skottsk, 4...exd4 5.Nxd4 Bb4
C47.28=Fyra Springare: Skottsk, 4...exd4 5.Nxd4 Bb4 6.Nxc6 bxc6
C47.29=Fyra Springare: Skottsk, Huvudvarianten
C47.30=Fyra Springare: Skottsk, Huvudvarianten, 7...d5
C47.31=Fyra Springare: Skottsk, Huvudvarianten, 7...d5 8.exd5 cxd5
C47.32=Fyra Springare: Skottsk, Huvudvarianten, 8.exd5 cxd5 9.O-O O-O
C47.33=Fyra Springare: Skottsk, Huvudvarianten, 9.O-O O-O 10.Bg5 c6
C47.34=Fyra Springare: Skottsk, Huvudvarianten, 10.Bg5 c6 11.Na4
C47.35=Fyra Springare: Skottsk, Huvudvarianten, 10.Bg5 c6 11.Qf3
C47.36=Fyra Springare: Skottsk, Huvudvarianten, 10.Bg5 c6 11.Qf3 Be7
C48.1=Fyra Springare: Spanskt variant
C48.2=Fyra Springare: Spanskt, Rankenvarianten
C48.3=Fyra Springare: Spanskt, Spielmannvarianten
C48.4=Fyra Springare: Spanskt, 4...d6
C48.5=Fyra Springare: Spanskt, 4...d6 5.d4
C48.6=Fyra Springare: Spanskt, Klassiskt f�rsvar
C48.7=Fyra Springare: Spanskt, Klassiskt f�rsvar, 5.Nxe5
C48.8=Fyra Springare: Spanskt, Klassiskt f�rsvar, 5.O-O
C48.9=Fyra Springare: Spanskt, Klassisk, Bardelebenvarianten
C48.10=Fyra Springare: Spanskt, Klassisk, Marshallvarianten
C48.11=Fyra Springare: Rubinsteins motgambit
C48.12=Fyra Springare: Rubinstein, 5.Be2
C48.13=Fyra Springare: Rubinstein, 5.Nxe5
C48.14=Fyra Springare: Rubinstein, Bogoljubowvarianten
C48.15=Fyra Springare: Rubinstein, Hennebergervarianten
C48.16=Fyra Springare: Rubinstein, 5.Bc4
C48.17=Fyra Springare: Rubinstein, Avbytesvarianten
C48.18=Fyra Springare: Rubinstein, Avbytesvarianten
C48.19=Fyra Springare: Rubinstein, Avbytesvarianten, 8...Bc5
C48.20=Fyra Springare: Rubinstein, Avbytesvarianten, 8...Qe5+
C48.21=Fyra Springare: Rubinstein, 5.Ba4
C48.22=Fyra Springare: Rubinstein, 5.Ba4 Nxf3+
C48.23=Fyra Springare: Rubinstein, 5.Ba4 c6
C48.24=Fyra Springare: Rubinstein, 5.Ba4 c6 6.Nxe5
C48.25=Fyra Springare: Rubinstein, 5.Ba4 Bc5
C48.26=Fyra Springare: Rubinstein, 5.Ba4 Bc5 6.Nxe5
C49.1=Fyra Springare: 4.Bb5 Bb4
C49.2=Fyra Springare: 4.Bb5 Bb4 5.O-O
C49.3=Fyra Springare: 4.Bb5 Bb4 5.O-O O-O
C49.4=Fyra Springare: Gunsbergvarianten
C49.5=Fyra Springare: Nimzowitsch (Paulsen)varianten
C49.6=Fyra Springare: Dubbla l�pare, 6.d3
C49.7=Fyra Springare: Dubbla l�pare, 6.d3 Bxc3
C49.8=Fyra Springare: Janowski varianten
C49.9=Fyra Springare: Svenonius varianten
C49.10=Fyra Springare: Symmetriska varianten
C49.11=Fyra Springare: Symmetrisk, Maroczysystemet
C49.12=Fyra Springare: Symmetrisk, 7.Bg5
C49.13=Fyra Springare: Symmetrisk, Tarraschvarianten
C49.14=Fyra Springare: Symmetrisk, Pillsburyvarianten
C49.15=Fyra Springare: Symmetrisk, Blakevarianten
C49.16=Fyra Springare: Symmetrisk, 7.Bg5 Bxc3
C49.17=Fyra Springare: Symmetrisk, 7.Bg5 Bxc3
C49.18=Fyra Springare: Symmetrisk, 7.Bg5 Bxc3 8.bxc3 h6
C49.19=Fyra Springare: Symmetrisk, Metger frig�ra
C49.20=Fyra Springare: Symmetrisk, Metger, 10.d4
C49.21=Fyra Springare: Symmetrisk, Metger, Capablancavarianten
C49.22=Fyra Springare: Symmetrisk, Metger, 10.d4 Ne6
C49.23=Fyra Springare: Symmetrisk, Metger, 10.d4 Ne6 11.Bc1 Rd8
C49.24=Fyra Springare: Symmetrisk, Metger, 10.d4 Ne6 11.Bc1 c5
C50.1=Italienskt parti
C50.2=Italienskt: Rousseaus gambit
C50.3=Italienskt: Blackburne-Shillings gambit
C50.4=Italienskt: 3...d6
C50.5=Italienskt: Ungerskt f�rsvar
C50.6=Italienskt: Ungerskt f�rsvar, 4.d4 exd4
C50.7=Italienskt: Ungerskt f�rsvar, Tartakowervarianten
C50.8=Italienskt: Ungerskt f�rsvar, 4.d4 d6
C50.9=Giuoco Piano
C50.10=Giuoco Piano: Jeromes gambit
C50.11=Giuoco Piano: Rosentreters gambit
C50.12=Giuoco Piano: Trespringarvarianten
C50.13=Giuoco Piano: Fyrspringarvarianten
C50.14=Giuoco Piano: 4.O-O
C50.15=Giuoco Piano: 4.O-O Nf6
C50.16=Giuoco Piano: 4.O-O Nf6 5.Nc3
C50.17=Giuoco Pianissimo: 4.d3
C50.18=Giuoco Pianissimo: Lucchinis gambit
C50.19=Giuoco Pianissimo: Duboisvarianten
C50.20=Giuoco Pianissimo: 4.d3 Nf6
C50.21=Giuoco Pianissimo: 4.d3 Nf6 5.O-O
C50.22=Giuoco Pianissimo: 4.d3 Nf6 5.O-O d6
C50.23=Giuoco Pianissimo: Italienskt fyrspringar
C50.24=Giuoco Pianissimo: Italienskt fyrspringar, 5...d6
C50.25=Giuoco Pianissimo: Italienskt fyrspringar, 5...d6 6.Be3
C50.26=Giuoco Pianissimo: Canalvarianten
C50.27=Giuoco Pianissimo: Canal, 6...h6
C51.1=Evans gambit
C51.2=Avb�jd Evans gambit: 4...Be7
C51.3=Evans gambit: Heins motgambit
C51.4=Avb�jd Evans gambit
C51.5=Avb�jd Evans gambit, Cordelvarianten
C51.6=Avb�jd Evans gambit, 5.b5
C51.7=Avb�jd Evans gambit, Langevarianten
C51.8=Avb�jd Evans gambit, Pavlovvarianten
C51.9=Avb�jd Evans gambit, Hirschbachvarianten
C51.10=Avb�jd Evans gambit, Vasquezvarianten
C51.11=Avb�jd Evans gambit, Hickenvarianten
C51.12=Avb�jd Evans gambit, 5.a4
C51.13=Avb�jd Evans gambit, Showalter-varianten
C51.14=Antagen Evans gambit
C51.15=Antagen Evans gambit, 5.c3
C51.16=Evans gambit: Mayets f�rsvar
C51.17=Evans gambit: Stone-Wares f�rsvar
C51.18=Evans gambit: Anderssenvarianten
C51.19=Evans gambit: Anderssen, 6.Qb3
C51.20=Evans gambit: Anderssen, 6.d4
C51.21=Evans gambit: Cordelvarianten
C51.22=Evans gambit: Normalvarianten
C51.23=Evans gambit: Anderssenvarianten
C51.24=Evans gambit: Ulvestadvarianten
C51.25=Evans gambit: Paulsenvarianten
C51.26=Evans gambit: Morphyattack
C51.27=Evans gambit: G�ringattack
C51.28=Evans gambit: Steinitzvarianten
C51.29=Evans gambit: Normalvarianten
C51.30=Evans gambit: Fraserattack
C51.31=Evans gambit: Fraser-Mortimer attack
C52.1=Evans gambit: 5...Ba5
C52.2=Evans gambit: 5...Ba5 6.Qb3
C52.3=Evans gambit: 5...Ba5 6.O-O
C52.4=Evans gambit: 5...Ba5 6.O-O Nf6
C52.5=Evans gambit: Richardson-attack
C52.6=Evans gambit: 5...Ba5 6.O-O d6
C52.7=Evans gambit: 5...Ba5 6.O-O d6 7.d4
C52.8=Evans gambit: Waller-attack
C52.9=Evans gambit: Sanders-Alapinvarianten
C52.10=Evans gambit: Alapin-Steinitzvarianten
C52.11=Evans gambit: Laskers f�rsvar
C52.12=Evans gambit: 5...Ba5 6.d4
C52.13=Evans gambit: Leonhardtvarianten
C52.14=Evans gambit: 5...Ba5 6.d4 exd4
C52.15=Evans gambit: Kompromenterat f�rsvar
C52.16=Evans gambit: Kompromenterat f�rsvar, Paulsenvarianten
C52.17=Evans gambit: Kompromenterat f�rsvar, Pottervarianten
C52.18=Evans gambit: 5...Ba5 6.d4 d6
C52.19=Evans gambit: Sokolskyvarianten
C52.20=Evans gambit: Tartakower attack
C52.21=Evans gambit: Tartakower attack, 7...Qd7
C52.22=Evans gambit: Tartakower attack, 8.dxe5 Bb6
C52.23=Evans gambit: Tartakower attack, 8.dxe5 dxe5
C52.24=Evans gambit: Tartakower, Levenfishvarianten
C53.1=Giuoco Piano: 4.c3
C53.2=Giuoco Piano: La Bourdonnais-varianten
C53.3=Giuoco Piano: St�ngd variant
C53.4=Giuoco Piano: Centrum-kontrollvarianten
C53.5=Giuoco Piano: Tarraschvarianten
C53.6=Giuoco Piano: Mestelvarianten
C53.7=Giuoco Piano: Eisingervarianten
C54.1=Giuoco Piano: 4.c3 Nf6
C54.2=Giuoco Piano: Albins gambit
C54.3=Giuoco Piano: Birds attack
C54.4=Giuoco Piano: Birds attack
C54.5=Giuoco Pianissimo: 5.d3
C54.6=Giuoco Pianissimo: 5.d3 a6
C54.7=Giuoco Pianissimo: 5.d3 d6
C54.8=Giuoco Pianissimo: 5.d3 d6 6.Nbd2
C54.9=Giuoco Pianissimo: 5.d3 d6 6.O-O
C54.10=Giuoco Pianissimo: 5.d3 d6 6.O-O O-O
C54.11=Giuoco Piano: 5.d4
C54.12=Giuoco Piano: 6.e5
C54.13=Giuoco Piano: Ghulam Kassim-varianten
C54.14=Giuoco Piano: 6.e5 d5
C54.15=Giuoco Piano: Anderssenvarianten
C54.16=Giuoco Piano: 6.cxd4
C54.17=Giuoco Piano: 6.cxd4 Bb4+
C54.18=Giuoco Piano: Krakowvarianten
C54.19=Giuoco Piano: 6.cxd4 Bb4+ 7.Bd2
C54.20=Giuoco Piano: Krausevarianten
C54.21=Giuoco Piano: Greco attack
C54.22=Giuoco Piano: Greco attack
C54.23=Giuoco Piano: Bernsteinvarianten
C54.24=Giuoco Piano: Aitkenvarianten
C54.25=Giuoco Piano: Greco attack
C54.26=Giuoco Piano: Steinitzvarianten
C54.27=Giuoco Piano: M�ller (Therkatz) attack
C54.28=Giuoco Piano: M�ller-Herzogvarianten
C54.29=Giuoco Piano: M�ller, Barjonettattack
C55.1=Tv�springarf�rsvar
C55.2=Tv� springare: Deutz gambit
C55.3=Tv� springare: 4.O-O gambit, Rosentretervarianten
C55.4=Tv� springare: 4.O-O gambit, Holzhausen attack
C55.5=Tv� springare: 4.d3
C55.6=Tv� springare: 4.d3 h6
C55.7=Tv� springare: 4.d3 Be7
C55.8=Tv� springare: 4.d3 Be7 5.Bb3 O-O
C55.9=Tv� springare: 4.d3 Be7 5.c3
C55.10=Tv� springare: 4.d3 Be7 5.O-O
C55.11=Tv� springare: 4.d3 Be7 5.O-O O-O
C55.12=Tv� springare: 4.d3 Be7 5.O-O O-O 6.Bb3
C55.13=Tv� springare: 4.d3 Be7 5.O-O O-O 6.Bb3 d6 7.c3
C55.14=Tv� springare: 4.d3 Be7 5.O-O O-O 6.Re1
C55.15=Tv� springare: 4.d4
C55.16=Tv� springare: 4.d4 exd4
C55.17=Tv� springare: 4.d4 exd4 5.Nxd4
C55.18=Tv� springare: Perreuxvarianten
C55.19=Tv� springare: Modern variant
C55.20=Tv� springare: Modern, 5.e5 d5
C55.21=Tv� springare: Modern, Huvudvarianten
C55.22=Tv� springare: Modern, Huvudvarianten, 8.Bxc6 bxc6 9.O-O Bc5
C55.23=Tv� springare: 5.O-O
C55.24=Tv� springare: 5.O-O Be7
C55.25=Tv� springare: 5.O-O d6
C55.26=Tv� springare: Max Lange attack
C55.27=Tv� springare: Max Lange, Steinitzvarianten
C55.28=Tv� springare: Max Lange, Krausevarianten
C55.29=Tv� springare: Max Lange, 6.e5 d5
C55.30=Tv� springare: Max Lange, Schlechtervarianten
C55.31=Tv� springare: Max Lange, Bergervarianten
C55.32=Tv� springare: Max Lange, Marshallvarianten
C55.33=Tv� springare: Max Lange, Rubinsteinvarianten
C55.34=Tv� springare: Max Lange, Lomans f�rsvar
C56.1=Tv� springare: Klassisk
C56.2=Tv� springare: Klassisk, Nakhmansonvarianten
C56.3=Tv� springare: Klassisk, 6.Re1
C56.4=Tv� springare: Klassisk, 6.Re1 d5
C56.5=Tv� springare: Klassisk, Canalvarianten
C56.6=Tv� springare: Klassisk, 7.Bxd5
C56.7=Tv� springare: Klassisk, 7.Bxd5 Qxd5
C56.8=Tv� springare: Klassisk, 8.Nc3
C56.9=Tv� springare: Klassisk, 8.Nc3 Qd8
C56.10=Tv� springare: Klassisk, 8.Nc3 Qh5
C56.11=Tv� springare: Klassisk, 8.Nc3 Qh5 9.Nxe4 Be6 10.Bg5 Bd6
C56.12=Tv� springare: Klassisk, M�llervarianten
C56.13=Tv� springare: Klassisk, M�ller, 9.Nxe4
C56.14=Tv� springare: Klassisk, M�ller, 9.Nxe4 Be6
C56.15=Tv� springare: Klassisk, M�ller, 10.Bg5
C56.16=Tv� springare: Klassisk, Yurdansky attack
C56.17=Tv� springare: Klassisk, M�ller, 10.Neg5
C56.18=Tv� springare: Klassisk, M�ller, 10.Neg5 O-O-O 11.Nxe6 fxe6 12.Rxe6 Bd6
C56.19=Tv� springare: Klassisk, M�ller, 10.Bd2
C56.20=Tv� springare: Klassisk, M�ller, 10.Bd2 Qf5
C56.21=Tv� springare: Klassisk, M�ller, 10.Bd2 Qd5
C56.22=Tv� springare: Klassisk, M�ller, 10.Bd2 Bb4
C57.1=Tv� springare: 4.Ng5
C57.2=Tv� springare: Traxler (Wilkes-Barre)varianten
C57.3=Tv� springare: Traxler, 5.d4
C57.4=Tv� springare: Traxler, 5.Nxf7
C57.5=Tv� springare: Traxler, 5.Nxf7 & 6.Kxf2
C57.6=Tv� springare: Traxler, 5.Nxf7 & 6.Kf1
C57.7=Tv� springare: Traxler, 5.Nxf7 & 6.Kf1, Beyers 8...Bg4
C57.8=Tv� springare: Traxler, 5.Nxf7 & 6.Kf1, 8...Nd4
C57.9=Tv� springare: Traxler, 5.Nxf7 & 6.Kf1, Palkinvarianten
C57.10=Tv� springare: Traxler, 5.Nxf7 & 6.Kf1, Menovskyvarianten
C57.11=Tv� springare: Traxler, 5.Bxf7+
C57.12=Tv� springare: Traxler, 5.Bxf7+ Ke7 6.Bb3
C57.13=Tv� springare: Traxler, Chigorin/Pithartvarianten
C57.14=Tv� springare: 4.Ng5 d5
C57.15=Tv� springare: Klossvarianten
C57.16=Tv� springare: 4.Ng5 d5 5.exd5 Nxd5
C57.17=Tv� springare: Lolli attack
C57.18=Tv� springare: Lolli attack, Pinkusvarianten
C57.19=Tv� springare: Fegatello (Stekt Lever) attack
C57.20=Tv� springare: Fegatello, Leonhardtvarianten
C57.21=Tv� springare: Fegatello, Polerios f�rsvar
C57.22=Tv� springare: Ulvestadvarianten
C57.23=Tv� springare: Fritzvarianten
C57.24=Tv� springare: Fritzvarianten, Huvudvarianten
C57.25=Tv� springare: Fritz, 8.Nxf7
C57.26=Tv� springare: Fritz, 8.cxd5
C57.27=Tv� springare: Fritz, Paoli's 8.h4
C57.28=Tv� springare: Fritz, Grubervarianten (8.Ne4)
C57.29=Tv� springare: Fritz, Radchenkovarianten
C57.30=Tv� springare: Fritz, Berlinvarianten
C58.1=Tv� springare: Morphyvarianten (5...Na5)
C58.2=Tv� springare: Morphy, Kieseritskyvarianten
C58.3=Tv� springare: Morphy, Kieseritskyvarianten, 6...h6 7.Nf3 e4 8.Qe2
C58.4=Tv� springare: Morphy, Yankovichvarianten
C58.5=Tv� springare: Morphy, Maroczyvarianten
C58.6=Tv� springare: Morphy, Polerio (6.Bb5+)
C58.7=Tv� springare: Morphy, Polerio, 6...Bd7
C58.8=Tv� springare: Morphy, Polerio, 6...c6
C58.9=Tv� springare: Morphy, Bogoljubowvarianten
C58.10=Tv� springare: Morphy, Blackburnevarianten
C58.11=Tv� springare: Morphy, Paoli-varianten
C58.12=Tv� springare: Morphy, Colman-varianten
C58.13=Tv� springare: Morphy, 8.Be2
C59.1=Tv� springare: Morphy, 8.Be2 h6
C59.2=Tv� springare: Morphy, Steinitzvarianten
C59.3=Tv� springare: Morphy, Huvudvarianten 9.Nf3
C59.4=Tv� springare: Morphy, Huvudvarianten 9.Nf3 e4
C59.5=Tv� springare: Morphy, Huvudvarianten 9.Nf3 e4 10.Ne5
C59.6=Tv� springare: Morphy, Steinervarianten
C59.7=Tv� springare: Morphy, G�ringvarianten
C59.8=Tv� springare: Morphy, Gellervarianten
C59.9=Tv� springare: Huvudvarianten 10...Bd6
C59.10=Tv� springare: Huvudvarianten, 11.f4
C59.11=Tv� springare: Huvudvarianten, 11.f4 exf3
C59.12=Tv� springare: Huvudvarianten, 11.d4
C59.13=Tv� springare: Huvudvarianten, 11.d4 Qc7
C59.14=Tv� springare: Huvudvarianten, Knorrevarianten
C59.15=Tv� springare: Huvudvarianten, 11.d4 exd3
C59.16=Tv� springare: Huvudvarianten, 11.d4 exd3 12.Nxd3 Qc7
C59.17=Tv� springare: Huvudvarianten, 11.d4, Honfi-varianten
C60.1=Spanskt (Ruy Lopez)
C60.2=Spanskt: Spanskt motgambit
C60.3=Spanskt: 3...a5
C60.4=Spanskt: N�rnbergs variant
C60.5=Spanskt: Pollocks f�rsvar
C60.6=Spanskt: Lucenas f�rsvar
C60.7=Spanskt: Vinogradov-varianten
C60.8=Spanskt: Brentano-varianten
C60.9=Spanskt: Alapin-varianten
C60.10=Spanskt: Alapin, 4.c3
C60.11=Spanskt: Fianchetto (Smyslov) f�rsvar
C60.12=Spanskt: Fianchetto, 4.O-O
C60.13=Spanskt: Fianchetto, 4.d4
C60.14=Spanskt: Fianchetto, 4.d4 exd4 5.Bg5
C60.15=Spanskt: Fianchetto, 4.c3
C60.16=Spanskt: Cozios f�rsvar
C60.17=Spanskt: Cozio, 4.Nc3
C60.18=Spanskt: Cozio, Paulsen-varianten
C60.19=Spanskt: Cozio, 4.O-O
C60.20=Spanskt: Cozio, 4.O-O
C60.21=Spanskt: Cozio, 4.O-O g6
C60.22=Spanskt: Cozio, 4.O-O g6
C61.1=Spanskt: Birds f�rsvar
C61.2=Spanskt: Bird, 4.Bc4
C61.3=Spanskt: Bird, 4.Nxd4
C61.4=Spanskt: Bird, 4.Nxd4 exd4
C61.5=Spanskt: Bird, 5.d3
C61.6=Spanskt: Bird, 5.Bc4
C61.7=Spanskt: Bird, 5.O-O
C61.8=Spanskt: Bird, Paulsenvarianten
C61.9=Spanskt: Bird, 5.O-O c6
C61.10=Spanskt: Bird, 5.O-O c6 6.Bc4
C61.11=Spanskt: Bird, 5.O-O Bc5
C61.12=Spanskt: Bird, 5.O-O Bc5 6.d3
C61.13=Spanskt: Bird, 5.O-O Bc5 6.d3 c6
C61.14=Spanskt: Bird, 5.O-O Bc5 6.d3 c6 7.Bc4
C61.15=Spanskt: Bird, 5.O-O Bc5 6.d3 c6 7.Bc4 d5
C62.1=Spanskt: Gamla Steinitz
C62.2=Spanskt: Gamla Steinitz, 4.Bxc6+
C62.3=Spanskt: Gamla Steinitz, 4.O-O
C62.4=Spanskt: Gamla Steinitz, 4.c3
C62.5=Spanskt: Gamla Steinitz, 4.d4
C62.6=Spanskt: Gamla Steinitz, 4.d4 exd4
C62.7=Spanskt: Gamla Steinitz, 4.d4 exd4 5.Qxd4
C62.8=Spanskt: Gamla Steinitz, 4.d4 exd4 5.Nxd4
C62.9=Spanskt: Gamla Steinitz, 4.d4 Bd7
C62.10=Spanskt: Gamla Steinitz, 4.d4 Bd7 5.Nc3
C62.11=Spanskt: Gamla Steinitz, Nimzowitsch-attacken
C62.12=Spanskt: Gamla Steinitz, Semi-Durasvarianten
C63.1=Spanskt: Schliemann (J�nisch)
C63.2=Spanskt: Schliemann, 4.Qe2
C63.3=Spanskt: Schliemann, 4.exf5
C63.4=Spanskt: Schliemann, 4.d4
C63.5=Spanskt: Schliemann, 4.d3
C63.6=Spanskt: Schliemann, 4.d3 fxe4
C63.7=Spanskt: Schliemann, 4.d3 fxe4 5.dxe4 Nf6 6.O-O
C63.8=Spanskt: Schliemann, 4.Bxc6
C63.9=Spanskt: Schliemann, 4.Bxc6 dxc6
C63.10=Spanskt: Schliemann, 4.Nc3
C63.11=Spanskt: Schliemann, 4.Nc3 Nd4
C63.12=Spanskt: Schliemann, 4.Nc3 Nd4 5.Ba4
C63.13=Spanskt: Schliemann, 4.Nc3 Nf6
C63.14=Spanskt: Schliemann, 4.Nc3 Nf6 5.exf5
C63.15=Spanskt: Schliemann, 4.Nc3 fxe4
C63.16=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 Nf6
C63.17=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 Nf6 6.Qe2
C63.18=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 Nf6 6.Nxf6+
C63.19=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 d5
C63.20=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 d5 6.Nxe5
C63.21=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 d5 6.Nxe5 dxe4 7.Nxc6 Qd5
C63.22=Spanskt: Schliemann, 4.Nc3 fxe4 5.Nxe4 d5 6.Nxe5 dxe4 7.Nxc6 Qg5
C64.1=Spanskt: Klassisk f�rsvar
C64.2=Spanskt: Klassisk, Avbyte
C64.3=Spanskt: Klassisk, 4.c3
C64.4=Spanskt: Klassisk, Bodenvarianten
C64.5=Spanskt: Klassisk, Charousek-varianten
C64.6=Spanskt: Klassisk, 4.c3 Nge7
C64.7=Spanskt: Klassisk, 4.c3 Qf6
C64.8=Spanskt: Klassisk, Cordels gambit
C64.9=Spanskt: Klassisk, Cordels gambit, 5.d4
C64.10=Spanskt: Klassisk, 4.c3 Nf6
C64.11=Spanskt: Klassisk, 4.c3 Nf6 5.d4
C64.12=Spanskt: Klassisk, 4.c3 Nf6 5.d4 Bb6
C64.13=Spanskt: Klassisk, 4.O-O
C64.14=Spanskt: Klassisk, 4.O-O Nge7
C64.15=Spanskt: Klassisk, 4.O-O Qf6
C64.16=Spanskt: Klassisk, 4.O-O d6
C64.17=Spanskt: Klassisk, 4.O-O d6 5.c3
C64.18=Spanskt: Klassisk, 4.O-O Nd4
C64.19=Spanskt: Klassisk, Zaitsevvarianten
C64.20=Spanskt: Klassisk, 4.O-O Nd4 5.Bc4
C64.21=Spanskt: Klassisk, 4.O-O Nd4 5.Nxd4
C64.22=Spanskt: Klassisk, 4.O-O Nd4 5.Nxd4 Bxd4
C64.23=Spanskt: Klassisk, 4.O-O Nd4 5.Nxd4 Bxd4 6.c3
C64.24=Spanskt: Klassisk, 4.O-O Nd4 5.Nxd4 Bxd4 6.c3 Bb6
C64.25=Spanskt: Klassisk, 4.O-O Nd4 5.Nxd4 Bxd4 6.c3 Bb6 7.d4
C64.26=Spanskt: Klassisk, 6.c3 Bb6 7.d4 c6 8.Ba4
C64.27=Spanskt: Klassisk, 6.c3 Bb6 7.d4 c6 8.Ba4 d6 9.Na3
C65.1=Spanskt: Berlinf�rsvaret
C65.2=Spanskt: Berlin, 4.Qe2
C65.3=Spanskt: Berlin, 4.d4
C65.4=Spanskt: Berlin, 4.d4 exd4
C65.5=Spanskt: Berlin, Nyholms attack
C65.6=Spanskt: Berlin, 4.d3
C65.7=Spanskt: Berlin, Mortimervarianten
C65.8=Spanskt: Berlin, Mortimers f�lla
C65.9=Spanskt: Berlin, 4.d3 d6
C65.10=Spanskt: Berlin, Anderssenvarianten
C65.11=Spanskt: Berlin, Durasvarianten
C65.12=Spanskt: Berlin, 4.d3 d6 5.c3
C65.13=Spanskt: Berlin, 4.d3 Bc5
C65.14=Spanskt: Berlin, Kaufmannvarianten
C65.15=Spanskt: Berlin, 4.O-O
C65.16=Spanskt: Berlin, 4.O-O Be7
C65.17=Spanskt: Berlin, Beverwijkvarianten
C65.18=Spanskt: Berlin, Beverwijk, 5.c3
C65.19=Spanskt: Berlin, Beneluxvarianten
C65.20=Spanskt: Berlin, Beneluxvarianten, 7.Bg5
C65.21=Spanskt: Berlin, Beverwijk, 5.Nxe5
C66.1=Spanskt: St�ngt Berlin
C66.2=Spanskt: St�ngt Berlin, 5.d4
C66.3=Spanskt: St�ngt Berlin, Chigorinvarianten
C66.4=Spanskt: St�ngt Berlin, 5.d4 Bd7
C66.5=Spanskt: St�ngt Berlin, Wolfvarianten
C66.6=Spanskt: St�ngt Berlin, Hedgehog-varianten
C66.7=Spanskt: St�ngt Berlin, Tarraschs f�lla
C66.8=Spanskt: St�ngt Berlin, Bernsteinvarianten
C66.9=Spanskt: St�ngt Berlin, Showalter-varianten
C67.1=Spanskt: �ppet Berlin
C67.2=Spanskt: �ppet Berlin, 5.Qe2
C67.3=Spanskt: �ppet Berlin, 5.Re1
C67.4=Spanskt: �ppet Berlin, 5.Re1 Nd6 6.Nxe5
C67.5=Spanskt: �ppet Berlin, 5.d4
C67.6=Spanskt: �ppet Berlin, Rosenthalvarianten
C67.7=Spanskt: �ppet Berlin, 5...Be7
C67.8=Spanskt: Berlin, Minckwitzvarianten
C67.9=Spanskt: �ppet Berlin, 5...Be7 6.Qe2
C67.10=Spanskt: �ppet Berlin, Trifunovicvarianten
C67.11=Spanskt: �ppet Berlin, 5...Be7 6.Qd2 Nd6
C67.12=Spanskt: �ppet Berlin, Cordelvarianten
C67.13=Spanskt: �ppet Berlin, 5...Be7 6.Qd2 Nd6 7.Bxc6 bxc6 8.dxe5 Nb7
C67.14=Spanskt: �ppet Berlin, Pillsburyvarianten
C67.15=Spanskt: �ppet Berlin, Zukertortvarianten
C67.16=Spanskt: �ppet Berlin, Winawers attack
C67.17=Spanskt: �ppet Berlin, Huvudvarianten 9.Nc3 (Rio de Janerio)
C67.18=Spanskt: �ppet Berlin, 5.d4 Nd6
C67.19=Spanskt: �ppet Berlin, Showalter-varianten
C67.20=Spanskt: �ppet Berlin, 5.d4 Nd6 6.dxe5
C67.21=Spanskt: �ppet Berlin, 5.d4 Nd6 6.Bxc6
C67.22=Spanskt: �ppet Berlin, 5.d4 Nd6 6.Bxc6 dxc6
C67.23=Spanskt: �ppet Berlin, 5.d4 Nd6 6.Bxc6 dxc6 7.dxe5 Nf5
C67.24=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte
C67.25=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3
C67.26=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3 h6
C67.27=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3 Ke8
C67.28=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3 Ke8 10.Rd1
C67.29=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3 Ke8 10.h3
C67.30=Spanskt: �ppet Berlin, 5.d4 Nd6 Dambyte, 9.Nc3 Ke8 10.h3 a5
C68.1=Spanskt: 3...a6
C68.2=Spanskt: 3...a6 4.Bc4
C68.3=Spanskt: Avbytesvarianten
C68.4=Spanskt: Avbyte, 4...bxc6
C68.5=Spanskt: Avbyte, 4...dxc6
C68.6=Spanskt: Avbyte, Laskervarianten
C68.7=Spanskt: Avbyte, Alekhinevarianten
C68.8=Spanskt: Avbyte, Keresvarianten
C68.9=Spanskt: Avbyte, Keres, 5...f6
C68.10=Spanskt: Avbyte, Romanovskyvarianten
C68.11=Spanskt: Avbyte, 5.Nc3 f6 6.d4
C68.12=Spanskt: Avbyte, 5.O-O
C68.13=Spanskt: Avbyte, 5.O-O Ne7
C68.14=Spanskt: Avbyte, 5.O-O Bd6
C68.15=Spanskt: Avbyte, 5.O-O Bd6 6.d4 exd4
C68.16=Spanskt: Avbyte, 5.O-O Bg4
C68.17=Spanskt: Avbyte, 5.O-O Bg4 6.h3
C68.18=Spanskt: Avbyte, Alapins gambit
C68.19=Spanskt: Avbyte, Alapins gambit, 7.d3 Qf6 8.Nbd2
C68.20=Spanskt: Avbyte, Bronsteinvarianten
C68.21=Spanskt: Avbyte, Bronstein, 6.d3
C68.22=Spanskt: Avbyte, Bronstein, 6.Na3
C68.23=Spanskt: Avbyte, Bronstein, 6.Na3 b5
C68.24=Spanskt: Avbyte, Bronstein, 6.Na3 Be6
C69.1=Spanskt: Avbyte, Gligoricvarianten
C69.2=Spanskt: Avbyte, Gligoric, 6.d4
C69.3=Spanskt: Avbyte, Gligoric, 6.d4 Bg4
C69.4=Spanskt: Avbyte, Gligoric, 6.d4 Bg4 7.c3
C69.5=Spanskt: Avbyte, Gligoric, 6.d4 Bg4 7.c3 Bd6
C69.6=Spanskt: Avbyte, Gligoric, 6.d4 Bg4 7.dxe5
C69.7=Spanskt: Avbyte, Gligoric, 6.d4 Bg4 Dambyte, 9.Rd3
C69.8=Spanskt: Avbyte, Gligoric, 6.d4 Bg4 Dambyte, 9.Rd3 Bd6
C69.9=Spanskt: Avbyte, Gligoric, 6.d4 exd4
C69.10=Spanskt: Avbyte, Gligoric, 6.d4 exd4 7.Qxd4
C69.11=Spanskt: Avbyte, Gligoric, 6.d4 exd4 7.Nxd4
C69.12=Spanskt: Avbyte, Gligoric, 6.d4 exd4 7.Nxd4 Ne7
C69.13=Spanskt: Avbyte, Gligoric, 6.d4 exd4 7.Nxd4 c5
C69.14=Spanskt: Avbyte, Gligoric, 8.Ne2
C69.15=Spanskt: Avbyte, Gligoric, 8.Nb3
C69.16=Spanskt: Avbyte, Gligoric, 8.Nb3 Dambyte
C69.17=Spanskt: Avbyte, Gligoric, 8.Nb3 Dambyte, 9...Bd7
C69.18=Spanskt: Avbyte, Gligoric, 8.Nb3 Dambyte, 9...Bg4
C69.19=Spanskt: Avbyte, Gligoric, 8.Nb3 Dambyte, 9...Bg4 10.f3 Be6
C70.1=Spanskt: 4.Ba4
C70.2=Spanskt: Brentanovarianten
C70.3=Spanskt: 4.Ba4 Be7
C70.4=Spanskt: Avb�jd Fianchetto
C70.5=Spanskt: Avb�jd Alapin
C70.6=Spanskt: Avb�jd Cozio
C70.7=Spanskt: Avb�jd Bird
C70.8=Spanskt: Avb�jd Klassisk
C70.9=Spanskt: Carovarianten
C70.10=Spanskt: Grazvarianten
C70.11=Spanskt: Taimanov (Kant)varianten
C70.12=Spanskt: Avb�jd Schliemann
C70.13=Spanskt: Avb�jd Schliemann, 5.d4
C70.14=Spanskt: Avb�jd Schliemann, 5.d4 exd4 6.e5
C71.1=Spanskt: Modern Steinitz f�rsvar
C71.2=Spanskt: Modern Steinitz, Trespringarvarianten
C71.3=Spanskt: Modern Steinitz, 5.d4
C71.4=Spanskt: Modern Steinitz, Noas Ark f�lla
C71.5=Spanskt: Modern Steinitz, Keresvarianten
C72.1=Spanskt: Modern Steinitz, 5.O-O
C72.2=Spanskt: Modern Steinitz, 5.O-O Ne7
C72.3=Spanskt: Modern Steinitz, 5.O-O Bg4
C72.4=Spanskt: Modern Steinitz, 5.O-O Bg4 6.h3
C72.5=Spanskt: Modern Steinitz, 5.O-O Bd7
C72.6=Spanskt: Modern Steinitz, 5.O-O Bd7 6.d4
C73.1=Spanskt: Modern Steinitz, Richtervarianten
C73.2=Spanskt: Modern Steinitz, Richtervarianten
C73.3=Spanskt: Modern Steinitz, Richtervarianten
C73.4=Spanskt: Modern Steinitz, Alapinvarianten
C74.1=Spanskt: Modern Steinitz, 5.c3
C74.2=Spanskt: Modern Steinitz, 5.c3 g6
C74.3=Spanskt: Modern Steinitz, Siestavarianten
C74.4=Spanskt: Modern Steinitz, Siesta, 6.exf5
C74.5=Spanskt: Modern Steinitz, Siesta, Kopayevvarianten
C74.6=Spanskt: Modern Steinitz, Siesta, Kopayev, Huvudvarianten
C75.1=Spanskt: Modern Steinitz, 5.c3 Bd7
C75.2=Spanskt: Modern Steinitz, 5.c3 Bd7 6.O-O
C75.3=Spanskt: Modern Steinitz, 5.c3 Bd7 6.d4
C75.4=Spanskt: Modern Steinitz, 5.c3 Bd7 6.d4 Nf6
C75.5=Spanskt: Modern Steinitz, Rubinsteinvarianten
C75.6=Spanskt: Modern Steinitz, Rubinstein, 7.Bb3
C75.7=Spanskt: Modern Steinitz, Rubinstein, 7.Be3
C76.1=Spanskt: Modern Steinitz, Bronsteinvarianten
C76.2=Spanskt: Modern Steinitz, Bronstein, 7.O-O
C76.3=Spanskt: Modern Steinitz, Bronstein, 7.O-O Bg7 8.Re1
C76.4=Spanskt: Modern Steinitz, Bronstein, 7.O-O Bg7 8.dxe5
C76.5=Spanskt: Modern Steinitz, Bronstein, 7.O-O Bg7 8.dxe5 dxe5
C76.6=Spanskt: Modern Steinitz, Bronstein, 7.O-O Bg7 8.dxe5 Nxe5
C76.7=Spanskt: Modern Steinitz, Bronstein, 7.O-O Bg7 8.d5
C77.1=Spanskt: Morphys f�rsvar
C77.2=Spanskt: Anderssenvarianten
C77.3=Spanskt: Anderssen, 5...b5
C77.4=Spanskt: Anderssen, 5...d6
C77.5=Spanskt: Durasvarianten
C77.6=Spanskt: Anderssen, 5...d6 6.c3
C77.7=Spanskt: Anderssen, 5...d6 6.c3 g6
C77.8=Spanskt: Fyrspringar (Tarrasch)varianten
C77.9=Spanskt: Avb�jt Avbyte
C77.10=Spanskt: Centrumattack
C77.11=Spanskt: Centrumattack, 5...b5
C77.12=Spanskt: Centrumattack, 5...Nxd4
C77.13=Spanskt: Centrumattack, 5...Nxe4
C77.14=Spanskt: Centrumattack, 5...Be7
C77.15=Spanskt: Centrumattack, 5...exd4
C77.16=Spanskt: Wormalds attack
C77.17=Spanskt: Wormalds attack, 5...Be7
C77.18=Spanskt: Wormalds attack, 5...b5
C77.19=Spanskt: Wormalds attack, 5...b5 6.Bb3 Bc5
C77.20=Spanskt: Wormalds attack, 5...b5 6.Bb3 Bc5 7.c3
C77.21=Spanskt: Wormalds attack, 5...b5 6.Bb3 Be7
C77.22=Spanskt: Wormalds attack, Gr�nfeldvarianten
C78.1=Spanskt: 5.O-O
C78.2=Spanskt: M�llers f�rsvar
C78.3=Spanskt: M�llers f�rsvar, 6.Nxe5
C78.4=Spanskt: M�llers f�rsvar, 6.c3
C78.5=Spanskt: 5.O-O b5
C78.6=Spanskt: 5.O-O b5 6.Bb3
C78.7=Spanskt: 5.O-O b5 6.Bb3 d6
C78.8=Spanskt: Rabinovich-varianten
C78.9=Spanskt: 5.O-O b5 6.Bb3 Be7
C78.10=Spanskt: 5.O-O b5 6.Bb3 Be7
C78.11=Spanskt: 5.O-O b5 6.Bb3 Bc5
C78.12=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.Nxe5
C78.13=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.Nxe5
C78.14=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.c3
C78.15=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.c3 d6
C78.16=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.c3 d6 8.d4
C78.17=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.a4
C78.18=Spanskt: 5.O-O b5 6.Bb3 Bc5 7.a4 Rb8
C78.19=Spanskt: Archangelsk-varianten
C78.20=Spanskt: Archangelsk, 7.d4
C78.21=Spanskt: Archangelsk, 7.d3
C78.22=Spanskt: Archangelsk, 7.d3 Be7
C78.23=Spanskt: Archangelsk, 7.c3
C78.24=Spanskt: Archangelsk, 7.c3 Nxe4
C78.25=Spanskt: Archangelsk, 7.Re1
C78.26=Spanskt: Archangelsk, 7.Re1 Bc5
C78.27=Spanskt: Archangelsk, 7.Re1 Bc5 8.c3 d6
C78.28=Spanskt: Archangelsk, Huvudvarianten
C78.29=Spanskt: Archangelsk, Huvudvarianten, 10.a4
C78.30=Spanskt: Archangelsk, Huvudvarianten, 10.Bg5
C78.31=Spanskt: Archangelsk, Huvudvarianten, 10.Be3
C79.1=Spanskt: Avb�jd Steinitz
C79.2=Spanskt: Avb�jd Steinitz, 6.c3
C79.3=Spanskt: Avb�jd Steinitz, 6.Re1
C79.4=Spanskt: Avb�jd Steinitz, Avbyte
C79.5=Spanskt: Avb�jd Steinitz, Lipnitskyvarianten
C79.6=Spanskt: Avb�jd Steinitz, Rubinsteinvarianten
C79.7=Spanskt: Avb�jd Steinitz, BoleSlavisksky-varianten
C80.1=Spanskt: �ppet
C80.2=Spanskt: �ppet, Knorrevarianten
C80.3=Spanskt: �ppet, Tartakowervarianten
C80.4=Spanskt: �ppet, 6.Re1
C80.5=Spanskt: �ppet, 6.Re1 Nc5 7.Bxc6
C80.6=Spanskt: �ppet, 6.d4
C80.7=Spanskt: �ppet, Rigavarianten
C80.8=Spanskt: �ppet, 6.d4 Be7
C80.9=Spanskt: �ppet, 6.d4 b5
C80.10=Spanskt: �ppet, Friess attack
C80.11=Spanskt: �ppet, Richtervarianten
C80.12=Spanskt: �ppet, 7.Bb3
C80.13=Spanskt: �ppet, 7.Bb3 d5
C80.14=Spanskt: �ppet, 7.Bb3 d5 8.a4
C80.15=Spanskt: �ppet, Schlechters f�rsvar
C80.16=Spanskt: �ppet, Schlecter, Bergervarianten
C80.17=Spanskt: �ppet, Harksens gambit
C80.18=Spanskt: �ppet, 8.Nxe5
C80.19=Spanskt: �ppet, 8.dxe5
C80.20=Spanskt: �ppet, Zukertortvarianten
C80.21=Spanskt: �ppet, 8...Be6
C80.22=Spanskt: �ppet, 8...Be6 9.a4
C80.23=Spanskt: �ppet, 8...Be6 9.Be3
C80.24=Spanskt: �ppet, Bernsteinvarianten
C80.25=Spanskt: �ppet, Bernstein, 9...Bc5
C80.26=Spanskt: �ppet, Bernstein, 9...Nc5
C80.27=Spanskt: �ppet, Bernstein, 9...Nc5 10.c3 d4
C80.28=Spanskt: �ppet, Bernstein, 11.cxd4
C80.29=Spanskt: �ppet, Bernstein, Karpovs gambit
C80.30=Spanskt: �ppet, Bernstein, 11.Bxe6
C81.1=Spanskt: �ppet, Keres attack
C81.2=Spanskt: �ppet, Keres attack, 9...Bc5
C81.3=Spanskt: �ppet, Keres attack, 9...Be7
C81.4=Spanskt: �ppet, Keres, Adamvarianten
C81.5=Spanskt: �ppet, Keres, 10.Rd1
C81.6=Spanskt: �ppet, Keres, 10.Rd1 O-O
C81.7=Spanskt: �ppet, Keres, 10.Rd1 O-O 11.c3
C81.8=Spanskt: �ppet, Keres, 10.Rd1 O-O 11.c4
C81.9=Spanskt: �ppet, Keres, 10.Rd1 O-O 11.c4 bxc4 12.Bxc4 Bc5
C81.10=Spanskt: �ppet, Keres, Ekstr�m-varianten
C82.1=Spanskt: �ppet, 9.c3
C82.2=Spanskt: �ppet, Berlinvarianten
C82.3=Spanskt: �ppet, Berlin, 10.Bc2
C82.4=Spanskt: �ppet, Berlin, 10.Bc2 Bg4
C82.5=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Re1
C82.6=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Nbd2
C82.7=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Nbd2 Be7
C82.8=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Nbd2 Be7 12.Re1
C82.9=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Nbd2 Be7 12.Re1 Qd7
C82.10=Spanskt: �ppet, Berlin, 10.Bc2 Bg4 11.Nbd2 Be7 12.Re1 O-O
C82.11=Spanskt: �ppet, Italiensk variant
C82.12=Spanskt: �ppet, Motzko attack
C82.13=Spanskt: �ppet, Motzko attack, Nenarokovvarianten
C82.14=Spanskt: �ppet, St. Petersburgvarianten
C82.15=Spanskt: �ppet, St. Petersburgvarianten
C82.16=Spanskt: �ppet, St. Petersburg, 11.Bc2
C82.17=Spanskt: �ppet, St. Petersburg, 11.Bc2 f5
C82.18=Spanskt: �ppet, Baguiovarianten
C82.19=Spanskt: �ppet, Baguio, 12.Nb3
C82.20=Spanskt: �ppet, Dilworthvarianten
C82.21=Spanskt: �ppet, Dilworth, 12.Rxf2 f6 13.exf6
C82.22=Spanskt: �ppet, Dilworth, 14.Kxf2
C82.23=Spanskt: �ppet, Dilworth, 14.Kxf2 Qxf6 15.Nf1
C82.24=Spanskt: �ppet, Dilworth, 14.Kxf2 Qxf6 15.Kg1
C82.25=Spanskt: �ppet, Dilworth, 14.Kxf2 Qxf6 15.Kg1 g5
C83.1=Spanskt: �ppet, Klassiskt f�rsvar
C83.2=Spanskt: �ppet, Klassisk, 10.Re1
C83.3=Spanskt: �ppet, Klassisk, Tarrasch Trap
C83.4=Spanskt: �ppet, Klassisk, Breslauvarianten
C83.5=Spanskt: �ppet, Klassisk, 10.Be3
C83.6=Spanskt: �ppet, Klassisk, 10.Nbd2
C83.7=Spanskt: �ppet, Klassisk, 10.Nbd2 Nc5
C83.8=Spanskt: �ppet, Klassisk, 10.Nbd2 O-O
C83.9=Spanskt: �ppet, Klassisk, Malkinvarianten
C83.10=Spanskt: �ppet, Klassisk, 10.Nbd2 O-O 11.Bc2
C83.11=Spanskt: �ppet, Klassisk, 10.Nbd2 O-O 11.Bc2 f5 12.exf6
C83.12=Spanskt: �ppet, Klassisk, 10.Nbd2 O-O 11.Bc2 f5 12.Nb3
C84.1=Spanskt: St�ngt system
C84.2=Spanskt: St�ngt, 6.Nc3
C84.3=Spanskt: St�ngt, 6.Nc3 b5
C84.4=Spanskt: St�ngt, 6.Nc3 b5 7.Bb3
C84.5=Spanskt: St�ngt, 6.Nc3 b5 7.Bb3 d6
C84.6=Spanskt: St�ngt, 6.Nc3 b5 7.Bb3 d6 8.Nd5
C84.7=Spanskt: St�ngt, 6.d3
C84.8=Spanskt: St�ngt, 6.d3 b5
C84.9=Spanskt: St�ngt, 6.d3 b5
C84.10=Spanskt: St�ngt, Centrumattack
C84.11=Spanskt: St�ngt, Centrumattack
C84.12=Spanskt: St�ngt, Centrumattack, 7.e5
C84.13=Spanskt: St�ngt, Centrumattack, 7.e5 Ne4
C84.14=Spanskt: St�ngt, Centrumattack, Baskisk gambit
C84.15=Spanskt: St�ngt, Centrumattack, Antagen baskisk gambit
C84.16=Spanskt: St�ngt, Centrumattack, 7.e5 Ne4 8.b4
C84.17=Spanskt: St�ngt, Centrumattack, 7.e5 Ne4 8.Nxd4
C84.18=Spanskt: St�ngt, Centrumattack, 7.e5 Ne4 8.Nxd4 Nxd4
C84.19=Spanskt: St�ngt, Centrumattack, 7.e5 Ne4 8.Nxd4 O-O
C84.20=Spanskt: St�ngt, Centrumattack, 7.Re1
C84.21=Spanskt: St�ngt, Centrumattack, 7.Re1 b5
C84.22=Spanskt: St�ngt, Centrumattack, 7.Re1 b5 8.e5
C84.23=Spanskt: St�ngt, Centrumattack, 7.Re1 b5 8.e5 Nxe5
C84.24=Spanskt: St�ngt, Centrumattack, 7.Re1 b5 8.e5 Nxe5 9.Rxe5
C84.25=Spanskt: St�ngt, Centrumattack, 7.Re1 O-O
C84.26=Spanskt: St�ngt, Centrumattack, 7.Re1 O-O 8.e5 Ne8
C84.27=Spanskt: St�ngt, Centrumattack, 7.Re1 O-O 8.e5 Ne8 9.c3
C84.28=Spanskt: St�ngt, Centrumattack, 7.Re1 O-O 8.e5 Ne8 9.Bf4
C85.1=Spanskt: St�ngt, Avbyte
C85.2=Spanskt: St�ngt, Avbyte
C85.3=Spanskt: St�ngt, Avbyte, 7.Qe2
C85.4=Spanskt: St�ngt, Avbyte, 7.Qe1
C85.5=Spanskt: St�ngt, Avbyte, 7.Qe1 Nd7
C85.6=Spanskt: St�ngt, Avbyte, 7.Qe1 Nd7 8.b3
C85.7=Spanskt: St�ngt, Avbyte, 7.d3
C85.8=Spanskt: St�ngt, Avbyte, 7.d3 Nd7
C85.9=Spanskt: St�ngt, Avbyte, 7.d3 Nd7 8.Nbd2
C85.10=Spanskt: St�ngt, Avbyte, 7.d3 Nd7 8.Nbd2 O-O 9.Nc4
C86.1=Spanskt: Worralls attack
C86.2=Spanskt: Worralls attack, 6...d6
C86.3=Spanskt: Worralls attack, 6...b5
C86.4=Spanskt: Worralls attack, 6...b5 7.Bb3
C86.5=Spanskt: Worralls attack, 7...d6
C86.6=Spanskt: Worralls attack, 7...d6 8.c3
C86.7=Spanskt: Worralls attack, 7...O-O
C86.8=Spanskt: Worralls attack, 7...O-O 8.a4
C86.9=Spanskt: Worralls attack, 7...O-O 8.c3
C86.10=Spanskt: Worralls attack, 7...O-O 8.c3 d6
C86.11=Spanskt: Worralls attack, 7...O-O 8.c3 d6 9.d4
C86.12=Spanskt: Worralls attack, 7...O-O 8.c3 d6 9.Rd1
C86.13=Spanskt: Worralls attack, 7...O-O 8.c3 d5
C86.14=Spanskt: Worralls attack, 7...O-O 8.c3 d5 9.exd5
C86.15=Spanskt: Worralls attack, 7...O-O 8.c3 d5 9.d3
C86.16=Spanskt: Worralls attack, 7...O-O 8.c3 d5 9.d3 Bb7
C87.1=Spanskt: St�ngt, 6.Re1
C87.2=Spanskt: St�ngt, Averbakh (Ryska) varianten
C87.3=Spanskt: St�ngt, Averbakh, 7.Bxc6+
C87.4=Spanskt: St�ngt, Averbakh, 7.c3
C87.9=Spanskt: St�ngt, Averbakh, 7.c3 Bg4
C87.10=Spanskt: St�ngt, Averbakh, 7.c3 Bg4 8.h3
C87.11=Spanskt: St�ngt, Averbakh, 7.c3 Bg4 8.d3
C87.5=Spanskt: St�ngt, Averbakh, 7.c3 O-O
C87.6=Spanskt: St�ngt, Averbakh, 7.c3 O-O 8.d4 Bd7
C87.7=Spanskt: St�ngt, Averbakh, 7.c3 O-O 8.d4 Bd7 9.Nbd2
C87.8=Spanskt: St�ngt, Averbakh, 7.c3 O-O 8.h3
C88.1=Spanskt: St�ngt, 6...b5
C88.2=Spanskt: St�ngt, 6...b5 7.Bb3
C88.3=Spanskt: St�ngt, Trajkovics motattack
C88.4=Spanskt: St�ngt 7...d6
C88.5=Spanskt: St�ngt, 7...d6 8.d4
C88.6=Spanskt: St�ngt, Noas Ark f�lla
C88.7=Spanskt: St�ngt 7...d6 8.c3
C88.8=Spanskt: St�ngt 7...d6 8.c3 Bg4
C88.9=Spanskt: St�ngt 7...d6 8.c3 Na5
C88.10=Spanskt: St�ngt, Leonhardtvarianten
C88.11=Spanskt: St�ngt, Ballavarianten
C88.12=Spanskt: St�ngt, 7...O-O
C88.13=Spanskt: St�ngt, 8.d3
C88.14=Spanskt: St�ngt, 8.d3 d6
C88.15=Spanskt: St�ngt, 8.h3
C88.16=Spanskt: St�ngt, 8.h3 Bb7 9.d3 d6
C88.17=Spanskt: St�ngt, Anti-Marshall 8.a4
C88.18=Spanskt: St�ngt, Anti-Marshall 8.a4 b4
C88.19=Spanskt: St�ngt, Anti-Marshall 8.a4 Bb7
C88.20=Spanskt: St�ngt, Anti-Marshall 8.a4 Bb7 9.d3
C88.21=Spanskt: St�ngt, Anti-Marshall 8.a4 Bb7 9.d3 d6
C88.22=Spanskt: St�ngt, Anti-Marshall 8.a4 Bb7 9.d3 d6 10.Nc3
C88.23=Spanskt: St�ngt, Anti-Marshall 8.a4 Bb7 9.d3 d6 10.c3
C88.24=Spanskt: St�ngt, 8.c3
C89.1=Spanskt: Marshalls motattack
C89.2=Spanskt: Marshall, 9.exd5
C89.3=Spanskt: Marshall, Herman, Steiner-varianten
C89.4=Spanskt: Marshall, 9.exd5 Nxd5
C89.5=Spanskt: Marshall, 9.exd5 Nxd5 10.Nxe5
C89.6=Spanskt: Marshall, 9.exd5 Nxd5 10.Nxe5 Nxe5
C89.7=Spanskt: Marshall, 11.Rxe5
C89.8=Spanskt: Marshall, 11.Rxe5 Nf6
C89.9=Spanskt: Marshall, 11.Rxe5 c6
C89.10=Spanskt: Marshall, 12.Bxd5
C89.11=Spanskt: Marshall, Kevitzvarianten
C89.12=Spanskt: Marshall, 12.d3
C89.13=Spanskt: Marshall, 12.d3 Bd6 13.Re1
C89.14=Spanskt: Marshall, 12.d3 Bd6 13.Re1 Qh4
C89.15=Spanskt: Marshall, Huvudvarianten (12.d4)
C89.16=Spanskt: Marshall, Huvudvarianten (12.d4 Bd6)
C89.17=Spanskt: Marshall, Huvudvarianten, 13.Re2
C89.18=Spanskt: Marshall, Huvudvarianten, 13.Re1
C89.19=Spanskt: Marshall, Huvudvarianten, 13.Re1 Qh4
C89.20=Spanskt: Marshall, Huvudvarianten, 13.Re1 Qh4 14.g3
C89.21=Spanskt: Marshall, Huvudvarianten, 14.g3 Qh3
C89.22=Spanskt: Marshall, Huvudvarianten, 15.Re4
C89.23=Spanskt: Marshall, Huvudvarianten, 15.Be3
C89.24=Spanskt: Marshall, Huvudvarianten, 15.Be3 Bg4
C89.25=Spanskt: Marshall, Huvudvarianten, 15.Be3 Bg4 16.Qd3
C89.26=Spanskt: Marshall, Huvudvarianten, 15.Be3 Bg4 16.Qd3 Rae8
C89.27=Spanskt: Marshall, Huvudvarianten, 16.Qd3 Rae8 17.Nd2
C89.28=Spanskt: Marshall, Huvudvarianten, Putta bonde-varianten
C89.29=Spanskt: Marshall, Huvudvarianten, Klassiska varianten
C89.30=Spanskt: Marshall, Huvudvarianten, Klassisk, 18.c4
C89.31=Spanskt: Marshall, Huvudvarianten, Klassisk, 18.Bxd5
C89.32=Spanskt: Marshall, Huvudvarianten, Klassisk, 18.Qf1
C89.33=Spanskt: Marshall, Huvudvarianten, Klassisk, 18.a4
C89.34=Spanskt: Marshall, Huvudvarianten, Klassisk, Spasskyvarianten
C89.35=Spanskt: Marshall, Huvudvarianten, Klassisk, 18.a4 f5
C90.1=Spanskt: St�ngt, 8...d6
C90.2=Spanskt: St�ngt, Lutikovvarianten
C90.3=Spanskt: St�ngt, Suetinvarianten
C90.4=Spanskt: St�ngt, 8...d6 9.a4
C90.5=Spanskt: St�ngt, 8...d6 9.a4 Bg4
C90.6=Spanskt: St�ngt, Pilnikvarianten
C90.7=Spanskt: St�ngt, Pilnik, 9...h6
C90.8=Spanskt: St�ngt, Pilnik, 9...Na5
C90.9=Spanskt: St�ngt, Pilnik, 9...Na5
C90.10=Spanskt: St�ngt, Pilnik, 9...Na5
C90.11=Spanskt: St�ngt, Pilnik, 11.Nbd2
C90.12=Spanskt: St�ngt, Pilnik, 11.Nbd2 Qc7
C90.13=Spanskt: St�ngt, Pilnik, 11.Nbd2 Nc6
C90.14=Spanskt: St�ngt, Pilnik, 11.Nbd2 Re8
C90.15=Spanskt: St�ngt, Pilnik, 12.Nf1
C90.16=Spanskt: St�ngt, Pilnik, 12.Nf1 Nc6
C90.17=Spanskt: St�ngt, Pilnik, 12.Nf1 Bf8
C90.18=Spanskt: St�ngt, Pilnik, 12.Nf1 h6
C91.1=Spanskt: St�ngt, 9.d4
C91.2=Spanskt: St�ngt, Bogoljubowvarianten
C91.3=Spanskt: St�ngt, Bogoljubow, 10.Be3
C91.4=Spanskt: St�ngt, Bogoljubow, 10.Be3 exd4
C91.5=Spanskt: St�ngt, Bogoljubow, 10.d5
C91.6=Spanskt: St�ngt, Bogoljubow, 10.d5 Na5
C91.7=Spanskt: St�ngt, Bogoljubow, 10.d5 Na5
C91.8=Spanskt: St�ngt, Bogoljubow, 10.d5 Na5 11.Bc2 Qc8
C91.9=Spanskt: St�ngt, Bogoljubow, 10.d5 Na5 11.Bc2 c6
C91.10=Spanskt: St�ngt, Bogoljubow, 10.d5 Na5 11.Bc2 c6 12.h3 Bc8
C92.1=Spanskt: St�ngt, 9.h3
C92.2=Spanskt: St�ngt, Keresvarianten
C92.3=Spanskt: St�ngt, Kholmovvarianten
C92.4=Spanskt: St�ngt, Kholmov, 11.Qxb3
C92.5=Spanskt: St�ngt, Karpovvarianten
C92.6=Spanskt: St�ngt, Karpovvarianten, 10.d4 Bf6
C92.7=Spanskt: St�ngt, Karpovvarianten, 10.d4 Bf6 11.a4
C92.8=Spanskt: St�ngt, Karpovvarianten, 10.d4 Bf6 11.a4 Bb7 12.Na3
C92.9=Spanskt: St�ngt, Zaitsev (Flohr)varianten
C92.10=Spanskt: St�ngt, Zaitsev, 10.d4
C92.11=Spanskt: St�ngt, Zaitsev, 10.d4 Re8
C92.12=Spanskt: St�ngt, Zaitsev, 11.Ng5
C92.13=Spanskt: St�ngt, Zaitsev, 11.Nbd2
C92.14=Spanskt: St�ngt, Zaitsev, 11.Nbd2 Bf8 12.d5 Nb8
C92.15=Spanskt: St�ngt, Zaitsev, 12.Bc2
C92.16=Spanskt: St�ngt, Zaitsev, 12.a3
C92.17=Spanskt: St�ngt, Zaitsev, 12.a4
C92.18=Spanskt: St�ngt, Zaitsev, 12.a4 h6
C92.19=Spanskt: St�ngt, Zaitsev, 12.a4 h6 13.Bc2
C92.20=Spanskt: St�ngt, Zaitsev, 12.a4 h6 13.Bc2 exd4
C92.21=Spanskt: St�ngt, Zaitsev, 12.a4 h6 13.Bc2 exd4 14.cxd4 Nb4 15.Bb1 c5
C93.1=Spanskt: St�ngt, Smyslovs f�rsvar
C93.2=Spanskt: St�ngt, Smyslov, 10.d4 Re8
C93.3=Spanskt: St�ngt, Smyslov, 10.d4 Re8 11.a4
C93.4=Spanskt: St�ngt, Smyslov, 10.d4 Re8 11.Be3
C93.5=Spanskt: St�ngt, Smyslov, 10.d4 Re8 11.Nbd2
C93.6=Spanskt: St�ngt, Smyslov, 10.d4 Re8 11.Nbd2 Bf8
C93.7=Spanskt: St�ngt, Smyslov, 12.a3
C93.8=Spanskt: St�ngt, Smyslov, 12.Bc2
C93.9=Spanskt: St�ngt, Smyslov, 12.Nf1
C93.10=Spanskt: St�ngt, Smyslov, 12.Nf1 Bb7
C93.11=Spanskt: St�ngt, Smyslov, 12.Nf1 Bd7
C94.1=Spanskt: St�ngt, Breyer f�rsvar
C94.2=Spanskt: St�ngt, Breyer, Matulovicvarianten
C94.3=Spanskt: St�ngt, Breyer, 10.d3
C94.4=Spanskt: St�ngt, Breyer, 10.d3 Nbd7
C94.5=Spanskt: St�ngt, Breyer, 10.d3 Nbd7 11.Nbd2
C94.6=Spanskt: St�ngt, Breyer, 10.d3 Nbd7 11.Nbd2 Bb7
C95.1=Spanskt: St�ngt, Breyer, 10.d4
C95.2=Spanskt: St�ngt, Breyer, 10.d4 Bb7
C95.3=Spanskt: St�ngt, Breyer, 10.d4 Nbd7
C95.4=Spanskt: St�ngt, Breyer, Simaginvarianten
C95.5=Spanskt: St�ngt, Breyer, 10.d4 Nbd7 11.Bg5
C95.6=Spanskt: St�ngt, Breyer, Arsenievvarianten
C95.7=Spanskt: St�ngt, Breyer, Arseniev, 11...c6
C95.8=Spanskt: St�ngt, Breyer, 10.d4 Nbd7 11.Nbd2
C95.9=Spanskt: St�ngt, Breyer, 10.d4 Nbd7 11.Nbd2 Bb7
C95.10=Spanskt: St�ngt, Breyer, 10.d4 Nbd7 11.Nbd2 Bb7 12.a4
C95.11=Spanskt: St�ngt, Breyer, 10.d4 Nbd7 11.Nbd2 Bb7 12.Bc2
C95.12=Spanskt: St�ngt, Breyer, Gligoricvarianten
C95.13=Spanskt: St�ngt, Breyer, Huvudvarianten
C95.14=Spanskt: St�ngt, Breyer, Huvudvarianten, 13.b4
C95.15=Spanskt: St�ngt, Breyer, Huvudvarianten, 13.a4
C95.16=Spanskt: St�ngt, Breyer, Huvudvarianten, 13.Nf1
C95.17=Spanskt: St�ngt, Breyer, Huvudvarianten, 13.Nf1 Bf8
C95.18=Spanskt: St�ngt, Breyer, Huvudvarianten, 13.Nf1 Bf8 14.Ng3
C95.19=Spanskt: St�ngt, Breyer, Huvudvarianten, 14.Ng3 c5
C95.20=Spanskt: St�ngt, Breyer, Huvudvarianten, 14.Ng3 g6
C95.21=Spanskt: St�ngt, Breyer, Huvudvarianten, 14.Ng3 g6 15.b3
C95.22=Spanskt: St�ngt, Breyer, Huvudvarianten, 14.Ng3 g6 15.a4
C95.23=Spanskt: St�ngt, Breyer, Huvudvarianten, 15.a4 c5
C95.24=Spanskt: St�ngt, Breyer, Huvudvarianten, 15.a4 c5 16.d5 c4
C96.1=Spanskt: St�ngt, Chigorin
C96.2=Spanskt: St�ngt, Chigorin, 10.Bc2
C96.3=Spanskt: St�ngt, Chigorin, 10...c6
C96.4=Spanskt: St�ngt, Chigorin, Rossolimovarianten
C96.5=Spanskt: St�ngt, Chigorin, 10...Bb7
C96.6=Spanskt: St�ngt, Chigorin, 10...c5
C96.7=Spanskt: St�ngt, Chigorin, 11.d3
C96.8=Spanskt: St�ngt, Chigorin, 11.d3 Nc6
C96.9=Spanskt: St�ngt, Chigorin, 11.d4
C96.10=Spanskt: St�ngt, Chigorin, 11.d4 cxd4
C96.11=Spanskt: St�ngt, Chigorin, 11.d4 Bb7
C96.12=Spanskt: St�ngt, Chigorin, 11.d4 Bb7 12.Nbd2
C96.13=Spanskt: St�ngt, Chigorin, Borisenkovarianten
C96.14=Spanskt: St�ngt, Chigorin, Keresvarianten
C96.15=Spanskt: St�ngt, Chigorin, Keres, 11.Nbd2 cxd4
C97.1=Spanskt: St�ngt, Chigorin, 11.d4 Qc7
C97.2=Spanskt: St�ngt, Chigorin, 11.d4 Qc7 12.d5
C97.3=Spanskt: St�ngt, Chigorin, 11.d4 Qc7 12.d5 c4
C97.4=Spanskt: St�ngt, Chigorin, 11.d4 Qc7 12.Nbd2
C97.5=Spanskt: St�ngt, Chigorin, 12...Bb7
C97.6=Spanskt: St�ngt, Chigorin, 12...Re8
C97.7=Spanskt: St�ngt, Chigorin, 12...Rd8
C97.8=Spanskt: St�ngt, Chigorin, 12...Bd7
C97.9=Spanskt: St�ngt, Chigorin, 12...Bd7 13.Nf1
C97.10=Spanskt: St�ngt, Chigorin, 12...Bd7 13.Nf1 Nc4
C97.11=Spanskt: St�ngt, Chigorin, 12...Bd7 13.Nf1 Rfe8
C97.12=Spanskt: St�ngt, Chigorin, Jugoslaviskt system
C98.1=Spanskt: St�ngt, Chigorin, 12...Nc6
C98.2=Spanskt: St�ngt, Chigorin, Rauzer attack
C98.3=Spanskt: St�ngt, Chigorin, Rauzer attack
C98.4=Spanskt: St�ngt, Chigorin, Rauzer, 14.Nf1
C98.5=Spanskt: St�ngt, Chigorin, Rauzer, 14.Nf1 Be6
C98.6=Spanskt: St�ngt, Chigorin, 12...Nc6 13.d5
C98.7=Spanskt: St�ngt, Chigorin, 12...Nc6 13.d5 Na5
C98.8=Spanskt: St�ngt, Chigorin, 12...Nc6 13.d5 Nd8
C98.9=Spanskt: St�ngt, Chigorin, 12...Nc6 13.d5 Nd8 14.Nf1
C98.10=Spanskt: St�ngt, Chigorin, 12...Nc6 13.d5 Nd8 14.a4
C99.1=Spanskt: St�ngt, Chigorin, 12...cxd4
C99.2=Spanskt: St�ngt, Chigorin, 12...cxd4 13.cxd4
C99.3=Spanskt: St�ngt, Chigorin, 13...Rd8
C99.4=Spanskt: St�ngt, Chigorin, 13...Bd7
C99.5=Spanskt: St�ngt, Chigorin, 13...Bd7 14.Nf1
C99.6=Spanskt: St�ngt, Chigorin, 13...Bd7 14.Nf1 Rac8 15.Ne3
C99.7=Spanskt: St�ngt, Chigorin, 13...Bb7
C99.8=Spanskt: St�ngt, Chigorin, 13...Bb7 14.Nf1
C99.9=Spanskt: St�ngt, Chigorin, 13...Bb7 14.Nf1 Rac8
C99.10=Spanskt: St�ngt, Chigorin, 13...Bb7 14.Nf1 Rac8 15.Re2
C99.11=Spanskt: St�ngt, Chigorin, 13...Bb7 14.d5
C99.12=Spanskt: St�ngt, Chigorin, 13...Bb7 14.d5 Rac8
C99.13=Spanskt: St�ngt, Chigorin, 13...Nc6
C99.14=Spanskt: St�ngt, Chigorin, 13...Nc6 14.a3
C99.15=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nf1
C99.16=Spanskt: St�ngt, Chigorin, 13...Nc6 14.d5
C99.17=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nb3
C99.18=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nb3 a5
C99.19=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nb3 a5 15.Be3 a4
C99.20=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nb3 a5 15.Be3 a4 16.Nbd2 Nb4
C99.21=Spanskt: St�ngt, Chigorin, 13...Nc6 14.Nb3 a5 15.Be3 a4 16.Nbd2 Bd7
D00.1=Dambondeparti
D00.2=Dambonde: 2.f4
D00.3=Dambonde: 2.g3
D00.4=Dambonde: 2.c3
D00.5=Dambonde: 2.c3 Nf6
D00.6=Dambonde: 2.c3 Nf6 3.Bf4
D00.7=Dambonde: 2.c3 Nf6 3.Bg5
D00.8=Dambonde: Masonvarianten
D00.9=Dambonde, Mason, Steinitz motgambit
D00.10=Dambonde: 2.e3
D00.11=Dambonde: 2.e3 Nf6
D00.12=Dambonde: Stonewallattack
D00.13=Hodgsonattack (Trompowsky vs. 1...d5)
D00.14=Hodgsonattack: Wellingvarianten
D00.15=Hodgsonattack: 2...f6
D00.16=Hodgsonattack: 2...g6
D00.17=Hodgsonattack: 2...c6
D00.18=Hodgsonattack, 2...h6
D00.19=Hodgsonattack: 2...h6 3.Bh4 c6
D00.20=Hodgsonattack: 2...h6 3.Bh4 c6 4.e3
D00.21=Hodgsonattack: 2...h6 3.Bh4 c6 4.e3 Qb6
D00.22=Trompowsky: 2...d5
D00.23=Trompowsky: 2...d5 3.Nd2
D00.24=Trompowsky: 2...d5 3.e3
D00.25=Trompowsky: 2...d5 3.e3 e6
D00.26=Trompowsky: 2...d5 3.Bxf6
D00.27=Trompowsky: 2...d5 3.Bxf6 gxf6
D00.28=Trompowsky: 2...d5 3.Bxf6 gxf6 4.e3
D00.29=Trompowsky: 2...d5 3.Bxf6 gxf6 4.e3 c5
D00.30=Trompowsky: 2...d5 3.Bxf6 exf6
D00.31=Trompowsky: 2...d5 3.Bxf6 exf6 4.e3
D00.32=Trompowsky: 2...d5 3.Bxf6 exf6 4.e3 Bf5
D00.33=Trompowsky: 2...d5 3.Bxf6 exf6 4.e3 c6
D00.34=Trompowsky: 2...d5 3.Bxf6 exf6 4.e3 Be6
D00.35=Trompowsky: 2...d5 3.Bxf6 exf6 4.e3 Bd6
D00.36=Blackmar-Diemers gambit (BDG): 2.e4
D00.37=Blackmar-Diemers: Beyers motgambit
D00.38=Blackmar-Diemers gambit (BDG): 2.e4 dxe4
D00.39=Blackmar-Diemers: T�lamodsgambit
D00.40=Blackmar-Diemers: Fritzattack
D00.41=Blackmar-Diemers: 2.e4 dxe4 3.Nc3
D00.42=Blackmar-Diemers: Grosshans f�rsvar
D00.43=Blackmar-Diemers: Zellers f�rsvar
D00.44=Blackmar-Diemers: Pohmlanns f�rsvar
D00.45=Blackmar-Diemers: Lembergers motgambit
D00.46=Blackmar-Diemers: Lembergers motgambit, Rassmussenattack
D00.47=Blackmar-Diemers: Lembergers motgambit, Sneiderattack
D00.48=Dambonde: Veresovattack
D00.49=Dambonde: Veresovattack
D00.50=Dambonde: Veresovattack
D00.51=Dambonde: Veresov, 3.Bf4
D00.52=Dambonde: Veresov, 3.Nf3
D00.53=Dambonde: Veresov, 3.Nf3 g6
D00.54=Dambonde: Anti-Kungsindisk
D00.55=Dambonde: Anti-Kungsindiskt, Huvudvarianten
D00.56=Blackmar-Diemers gambit (BDG)
D00.57=Blackmar-Diemers: Hubschs gambit
D00.58=Blackmar-Diemers: 3...dxe4
D00.59=Blackmar-Diemers: von Popiels attack
D00.60=Blackmar-Diemers: 4.f3
D00.61=Blackmar-Diemers: O'Kellys f�rsvar
D00.62=Blackmar-Diemers: Langeheineckes f�rsvar
D00.63=Blackmar-Diemers: Elberts motgambit
D00.64=Blackmar-Diemers: Weinspachs f�rsvar
D00.65=Blackmar-Diemers: Lambs f�rsvar
D00.66=Blackmar-Diemers: Vienna f�rsvar
D00.67=Blackmar-Diemers: Antagen
D00.68=Blackmar-Diemers: Ryders gambit
D00.69=Blackmar-Diemers: 4.f3 exf3 5.Nxf3
D00.70=Blackmar-Diemers: Gunderams f�rsvar
D00.71=Blackmar-Diemers: Tartakowers f�rsvar
D00.72=Blackmar-Diemers: Zieglers f�rsvar
D00.73=Blackmar-Diemers: Euwes f�rsvar
D00.74=Blackmar-Diemers: Bogoljubows f�rsvar
D01.1=Richter-Veresov attack
D01.2=Richter-Veresov: 3...Ne4
D01.3=Richter-Veresov: 3...e6
D01.4=Richter-Veresov: 3...h6
D01.5=Richter-Veresov: 3...g6
D01.6=Richter-Veresov: 3...c6
D01.7=Richter-Veresov: 3...c5
D01.8=Richter-Veresov: 3...Bf5
D01.9=Richter-Veresov: 3...Bf5 4.f3
D01.10=Richter-Veresov: 3...Bf5 4.Nf3
D01.11=Richter-Veresov: 3...Bf5 4.Bxf6
D01.12=Richter-Veresov: 3...Nbd7
D01.13=Richter-Veresov: 3...Nbd7 4.f3
D01.14=Richter-Veresov: 3...Nbd7 4.Nf3
D01.15=Richter-Veresov: 3...Nbd7 4.Nf3 h6
D01.16=Richter-Veresov: 3...Nbd7 4.Nf3 g6
D02.1=Dambonde: 2.Nf3
D02.2=Dambonde: 2.Nf3 g6
D02.3=Dambonde: 2.Nf3 Bg4
D02.4=Dambonde: 2.Nf3 c6
D02.5=Dambonde: London
D02.6=Dambonde: London, Alapinvarianten
D02.7=Dambonde: 2.Nf3 Bf5
D02.8=Dambonde: 2.Nf3 Bf5 3.e3
D02.9=Dambonde: 2.Nf3 Bf5 3.e3 c6
D02.10=Dambonde: 2.Nf3 Bf5 3.Bf4
D02.11=Dambonde: 2.Nf3 Bf5 3.Bf4 c6
D02.12=Dambonde: 2.Nf3 Bf5 3.Bf4 e6
D02.13=Dambonde: 2.Nf3 Nc6
D02.14=Dambonde: 2.Nf3 Nc6 3.Bf4
D02.15=Dambonde: 2.Nf3 Nc6 3.g3
D02.16=Dambonde: 2.Nf3 Nc6 3.g3 Bg4
D02.17=Dambonde: 2.Nf3 e6
D02.18=Dambonde: 2.Nf3 e6 3.g3
D02.19=Dambonde: 2.Nf3 e6 3.g3 c5
D02.20=Dambonde: 2.Nf3 e6 3.g3 c5
D02.21=Dambonde: 2.Nf3 e6 3.g3 c5
D02.22=Dambonde: 2.Nf3 e6 3.g3 c5
D02.23=Dambonde: Krausevarianten
D02.24=Dambonde: Krause, 3.c4
D02.25=Dambonde: Krause, Omv�nd slavisk
D02.26=Dambonde: Krause, Omv�nd avb�jd damgambit
D02.27=Dambonde: Krause, Omv�nd antagen damgambit
D02.28=Dambonde: 2.Nf3 Nf6
D02.29=Dambonde: 3.c3
D02.30=Dambonde: London
D02.31=Dambonde: London
D02.32=Dambonde: London
D02.33=Dambonde: London
D02.34=Dambonde: London
D02.35=Dambonde: London
D02.36=Dambonde: London
D02.37=Dambonde: 3.g3
D02.38=Dambonde: 3.g3 c6
D02.39=Dambonde: 3.g3 c6
D02.40=Dambonde: 3.g3 c6 4.Bg2 Bg4
D02.41=Dambonde: 3.g3 c6 4.Bg2 Bg4
D02.42=Dambonde: 3.g3 c6 4.Bg2 Bg4
D02.43=Dambonde: 3.g3 c6 4.Bg2 Bg4
D02.44=Dambonde: 3.g3 g6
D02.45=Dambonde: 3.g3 g6
D02.46=Dambonde: 3.g3 g6
A08.10=Retis: Antagen Kungsindisk, 2...c5 3.Bg2 Nc6 4.d4
D03.1=Torreattack (Tartakower)
D03.2=Torreattack: 3...Ne4
D03.3=Torreattack: 3...Ne4 4.Bf4
D03.4=Torreattack: 3...e6
D03.5=Torreattack: 3...e6 4.e3
D03.6=Torreattack: 3...e6 4.e3 Nbd7
D03.7=Torreattack: 3...e6 4.e3 Nbd7
D03.8=Torreattack: 3...e6 4.e3 c5
D03.9=Torreattack: 3...e6 4.e3 c5
D03.10=Torreattack: 3...e6 4.e3 c5
D03.11=Torreattack: 3...e6 4.e3 c5
D03.12=Torreattack: 3...g6
D03.13=Torreattack: 3...g6
D03.14=Torreattack: 3...g6
D03.15=Torreattack: 3...g6
D03.16=Torreattack: 3...g6 4.e3
D03.17=Torreattack: 3...g6 4.e3
D03.18=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2
D03.19=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O
D03.20=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.c3
D03.21=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.c3 Nbd7
D03.22=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.c3 Nbd7 7.Be2
D03.23=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.Bd3
D03.24=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.Bd3 c5
D03.25=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.Bd3 c5
D03.26=Torreattack: 3...g6 4.e3 Bg7 5.Nbd2 O-O 6.Bd3 c5 7.c3 Nbd7
D04.1=Dambonde: Colle
D04.2=Colle: 3...Bg4
D04.3=Colle: 3...Bf5
D04.4=Colle: 3...Bf5, Alekhinevarianten
D04.5=Colle: 3...g6
D04.6=Colle: 3...c6
D04.7=Colle: 3...c5
D04.8=Colle: 3...c5 4.c3
D04.9=Colle: 3...c5 4.c3 Nc6
D04.10=Colle: 3...c5 4.c3 Nbd7
D05.1=Colle: 3...e6
D05.2=Colle: 3...e6 4.Nbd2
D05.3=Colle: Zukertortvarianten
D05.4=Colle: 3...e6 4.Bd3
D05.5=Colle: Rubinsteins attack
D05.6=Colle: Rubinsteins attack, 5...Nc6
D05.7=Colle: 5.c3
D05.9=Colle: 5.c3 Nbd7
D05.8=Colle: 5.c3 Nc6
D06.1=Damgambit
D06.2=Avb�jd damgambit: �sterrikiskt f�rsvar
D06.3=Avb�jd damgambit: �sterrikiskt, Rubinsteinvarianten
D06.4=Avb�jd damgambit: �sterrikiskt, Rubinstein, 4.dxc5
D06.5=Avb�jd damgambit: �sterrikiskt, Rubinstein, 4.Nf3
D06.6=Avb�jd damgambit: �sterrikiskt, Rubinstein, 4.Nf3 cxd4
D06.7=Avb�jd damgambit: Marshalls f�rsvar
D06.8=Avb�jd damgambit: Marshalls f�rsvar, 3.Nc3
D06.9=Avb�jd damgambit: Marshalls f�rsvar, 3.Nf3
D06.10=Avb�jd damgambit: Marshalls f�rsvar, 3.cxd5
D06.11=Avb�jd damgambit: Marshalls f�rsvar, 3.cxd5 Nxd5
D06.12=Avb�jd damgambit: Marshalls f�rsvar, 3.cxd5 Nxd5 4.Nf3
D06.13=Avb�jd damgambit: Marshalls f�rsvar, 3.cxd5 Nxd5 4.e4
D06.14=Avb�jd damgambit: 2...Bf5
D06.15=Avb�jd damgambit: 2...Bf5 3.Qb3
D06.16=Avb�jd damgambit: 2...Bf5 3.Nc3
D06.17=Avb�jd damgambit: 2...Bf5 3.Nc3 e6
D06.18=Avb�jd damgambit: 2...Bf5 3.Nf3
D06.19=Avb�jd damgambit: 2...Bf5 3.Nf3 e6
D06.20=Avb�jd damgambit: 2...Bf5 3.Nf3 e6 4.Qb3
D06.21=Avb�jd damgambit: 2...Bf5 3.Nf3 e6 4.Nc3
D06.22=Avb�jd damgambit: 2...Bf5 3.Nf3 e6 4.Nc3 Nf6
D06.23=Avb�jd damgambit: 2...Bf5 3.cxd5
D06.24=Avb�jd damgambit: 2...Bf5 3.cxd5 Bxb1 4.Rxb1
D06.25=Avb�jd damgambit: 2...Bf5 3.cxd5 Bxb1 4.Qa4+
D06.26=Avb�jd damgambit: 2...Bf5 3.cxd5 Bxb1 4.Qa4+ c6 5.Rxb1
D07.1=Avb�jd damgambit: Chigorins f�rsvar
D07.2=Avb�jd damgambit: Chigorin, 3.cxd5
D07.3=Avb�jd damgambit: Chigorin, 3.cxd5, Huvudvarianten, 7.bxc3
D07.4=Avb�jd damgambit: Chigorin, 3.cxd5 Huvudvarianten, 7.Bxc3
D07.5=Avb�jd damgambit: Chigorin, 3.Nf3
D07.6=Avb�jd damgambit: Chigorin, Lazard gambit
D07.7=Avb�jd damgambit: Chigorin, 3.Nf3 Bg4
D07.8=Avb�jd damgambit: Chigorin, 3.Nf3 Bg4 4.Nc3
D07.9=Avb�jd damgambit: Chigorin, 3.Nf3 Bg4 4.cxd5
D07.10=Avb�jd damgambit: Chigorin, 3.Nf3 Bg4 4.cxd5 Bxf3 5.dxc6
D07.11=Avb�jd damgambit: Chigorin, 3.Nf3 Bg4 4.cxd5 Bxf3 5.gxf3
D07.12=Avb�jd damgambit: Chigorin, 3.Nc3
D07.13=Avb�jd damgambit: Chigorin, Tartakower gambit
D07.14=Avb�jd damgambit: Chigorin, 3.Nc3 Nf6
D07.15=Avb�jd damgambit: Chigorin, 3.Nc3 Nf6 4.Nf3
D07.16=Avb�jd damgambit: Chigorin, 3.Nc3 Nf6 4.Nf3 Bg4
D07.17=Avb�jd damgambit: Chigorin, 3.Nc3 dxc4
D07.18=Avb�jd damgambit: Chigorin, 3.Nc3 dxc4 4.d5
D07.19=Avb�jd damgambit: Chigorin, 3.Nc3 dxc4 4.Nf3
D07.20=Avb�jd damgambit: Chigorin, 3.Nc3 dxc4 4.Nf3 Nf6
D07.21=Avb�jd damgambit: Chigorin, 3.Nc3 dxc4 4.Nf3 Nf6 5.e4
D08.1=Avb�jd damgambit: Albins motgambit
D08.2=Avb�jd damgambit: Albin, 3.e3
D08.3=Avb�jd damgambit: Albin, 3.dxe5
D08.4=Avb�jd damgambit: Albin, 3.dxe5 d4
D08.5=Avb�jd damgambit: Albin, Laskers f�lla
D08.6=Avb�jd damgambit: Albin, 4.e4
D08.7=Avb�jd damgambit: Albin, 4.a3
D08.8=Avb�jd damgambit: Albin, 4.Nf3
D08.9=Avb�jd damgambit: Albin, 4.Nf3 Nc6
D08.10=Avb�jd damgambit: Albin, Alapinvarianten
D08.11=Avb�jd damgambit: Albin, Janowskivarianten
D08.12=Avb�jd damgambit: Albin, Baloghvarianten
D08.13=Avb�jd damgambit: Albin, Alapin, 5...Bg4
D08.14=Avb�jd damgambit: Albin, Krenoszvarianten
D08.15=Avb�jd damgambit: Albin, 4.Nf3 Nc6 5.a3
D08.16=Avb�jd damgambit: Albin, 4.Nf3 Nc6 5.a3 a5
D08.17=Avb�jd damgambit: Albin, 4.Nf3 Nc6 5.a3 Be6
D08.18=Avb�jd damgambit: Albin, 4.Nf3 Nc6 5.a3 Bg4
D08.19=Avb�jd damgambit: Albin, 4.Nf3 Nc6 5.a3 Bg4 6.Nbd2
D09.1=Avb�jd damgambit: Albin, 5.g3
D09.2=Avb�jd damgambit: Albin, 5.g3 Nge7
D09.3=Avb�jd damgambit: Albin, 5.g3 Bf5
D09.4=Avb�jd damgambit: Albin, 5.g3 Bg4
D09.5=Avb�jd damgambit: Albin, 5.g3 Bg4 6.Bg2 Qd7
D09.6=Avb�jd damgambit: Albin, 5.g3 Bg4 6.Bg2 Qd7 7.O-O O-O-O
D09.7=Avb�jd damgambit: Albin, 5.g3 Be6
D09.8=Avb�jd damgambit: Albin, 5.g3 Be6 6.b3
D09.9=Avb�jd damgambit: Albin, 5.g3 Be6 6.Bg2
D09.10=Avb�jd damgambit: Albin, 5.g3 Be6 6.Nbd2
D09.11=Avb�jd damgambit: Albin, 5.g3 Be6 6.Nbd2 Qd7
D09.12=Avb�jd damgambit: Albin, 5.g3 Be6 6.Nbd2 Qd7 7.Bg2
D09.13=Avb�jd damgambit: Albin, 5.g3 Be6 6.Nbd2 Qd7 7.Bg2 O-O-O
D09.14=Avb�jd damgambit: Albin, 5.g3 Be6 6.Nbd2 Qd7 7.Bg2 Nge7
D10.1=Slaviskt f�rsvar
D10.2=Diemer-Duhm gambit (DDG) mot Slavisk/Caro-Kann
D10.3=Slaviskt: 3.g3
D10.4=Slaviskt: 3.Bf4
D10.5=Slaviskt: Avbyte
D10.6=Slaviskt: Avbyte
D10.7=Slaviskt: Avbyte, 4.Bf4
D10.8=Slaviskt: Avbyte, 4.Nf3
D10.9=Slaviskt: Avbyte, 4.Nc3
D10.10=Slaviskt: Avbyte, 4.Nc3 Nf6
D10.11=Slaviskt: Avbyte, 4.Nc3 Nf6 5.Bf4
D10.12=Slaviskt: Avbyte, 4.Nc3 Nf6 5.Bf4 Nc6
D10.13=Slaviskt: Avbyte, 4.Nc3 Nf6 5.Bf4 Nc6 6.e3
D10.14=Slaviskt: Avbyte, 4.Nc3 Nf6 5.Bf4 Nc6 6.e3 a6
D10.15=Slaviskt: 3.e3
D10.16=Slaviskt: 3.e3 Bf5
D10.17=Slaviskt: 3.e3 Nf6
D10.18=Slaviskt: 3.Nc3
D10.19=Slaviskt: Winawers motgambit
D10.20=Slaviskt: Winawers motgambit, 4.cxd5
D10.21=Slaviskt: Winawers motgambit, 4.cxd5 cxd5 5.dxe5
D10.22=Slaviskt: Winawers motgambit, 4.cxd5 cxd5 5.Nf3
D10.23=Slaviskt: Antagen Winawers motgambit
D10.24=Slaviskt: Antagen Winawers motgambit, 6.Nd2
D10.25=Slaviskt: Antagen Winawers motgambit, 6.Bd2
D10.26=Slaviskt: 3.Nc3 dxc4
D10.27=Slaviskt: 3.Nc3 dxc4 4.a4
D10.28=Slaviskt: 3.Nc3 dxc4 4.e3
D10.29=Slaviskt: 3.Nc3 dxc4 4.e4
D10.30=Slaviskt: 3.Nc3 dxc4 4.e4 b5
D10.31=Slaviskt: 3.Nc3 dxc4 4.e4 b5 5.a4
D10.32=Slaviskt: 3.Nc3 Nf6
D10.33=Slaviskt: 3.Nc3 Nf6 4.Bg5
D10.34=Slaviskt: 3.Nc3 Nf6 4.Bg5 dxc4
D10.35=Slaviskt: 3.Nc3 Nf6 4.e3
D10.36=Slaviskt: 3.Nc3 Nf6 4.e3 Bf5
D10.37=Slaviskt: 3.Nc3 Nf6 4.e3 a6
D10.38=Slaviskt: 3.Nc3 Nf6 4.e3 a6 5.Bd3
D10.39=Slaviskt: 3.Nc3 Nf6 4.e3 a6 5.Qc2
D10.40=Slaviskt: 3.Nc3 Nf6 4.e3 a6 5.Qc2 b5
D11.1=Slaviskt: 3.Nf3
D11.2=Slaviskt: 3.Nf3 Bg4
D11.3=Slaviskt: 3.Nf3 Bf5
D11.4=Slaviskt: 3.Nf3 Bf5 4.Nc3
D11.5=Slaviskt: 3.Nf3 Bf5 4.Nc3 e6
D11.6=Slaviskt: 3.Nf3 Bf5 4.Nc3 e6 5.Qb3
D11.7=Slaviskt: 3.Nf3 dxc4
D11.8=Slaviskt: 3.Nf3 dxc4 4.Nc3
D11.9=Slaviskt: 3.Nf3 dxc4 4.e3
D11.10=Slaviskt: 3.Nf3 dxc4 4.e3 Be6
D11.11=Slaviskt: 3.Nf3 dxc4 4.e3 b5
D11.12=Slaviskt: 3.Nf3 dxc4 4.e3 b5 5.a4
D11.13=Slaviskt: 3.Nf3 dxc4 4.e3 b5 5.a4 e6
D11.14=Slaviskt: 3.Nf3 Nf6
D11.15=Slaviskt: 4.Qb3
D11.16=Slaviskt: 4.Qc2
D11.17=Slaviskt: 4.Qc2 g6 5.Bf4
D11.18=Slaviskt: Breyervarianten
D11.19=Slaviskt: Slaviskt-Reti system
D11.20=Slaviskt: Slaviskt-Reti system
D11.21=Slaviskt: Slaviskt-Reti system
D11.22=Slaviskt: Slaviskt-Reti system
D11.23=Slaviskt: Slaviskt-Reti system
D11.24=Slaviskt: Slaviskt-Reti system
D11.25=Slaviskt: Slaviskt-Reti system
D11.26=Slaviskt: Slaviskt-Reti system
D11.27=Slaviskt: Slaviskt-Reti system
D11.28=Slaviskt: Slavisk-Reti med b3
D11.29=Slaviskt: Slavisk-Reti med b3
D11.30=Slaviskt: Slavisk-Reti med b3
D11.31=Slaviskt: Slavisk-Reti med b3
D11.32=Slaviskt: Slavisk-Reti med b3
D11.33=Slaviskt: Slavisk-Reti med b3
D11.34=Slaviskt: Slavisk-Reti med b3
D11.35=Slaviskt: Slaviskt-Reti system
D11.36=Slaviskt: Slaviskt-Reti system
D11.37=Slaviskt: Slaviskt-Reti system
D11.38=Slaviskt: Slaviskt-Reti system
D11.39=Slaviskt: Slaviskt-Reti system
D11.40=Slaviskt: Slaviskt-Reti system
D11.41=Slaviskt: Slaviskt-Reti system
D11.42=Slaviskt: Slaviskt-Reti system
D11.43=Slaviskt: Slaviskt-Reti system
D11.44=Slaviskt: Slaviskt-Reti system
D11.45=Slaviskt: 4.e3
D11.46=Slaviskt: 4.e3 g6
D11.47=Slaviskt: 4.e3 a6
D11.48=Slaviskt: 4.e3 Bg4
D11.49=Slaviskt: 4.e3 Bg4
D12.1=Slaviskt: 4.e3 Bf5
D12.2=Slaviskt: 4.e3 Bf5 5.Qb3
D12.3=Slaviskt: 4.e3 Bf5 5.cxd5
D12.4=Slaviskt: 4.e3 Bf5 5.cxd5
D12.5=Slaviskt: 4.e3 Bf5 5.cxd5 cxd5 6.Qb3
D12.6=Slaviskt: 4.e3 Bf5 5.cxd5 cxd5 6.Qb3 Qc7
D12.7=Slaviskt: 4.e3 Bf5 5.cxd5 cxd5 6.Nc3
D12.8=Slaviskt: 4.e3 Bf5 5.cxd5 cxd5 6.Nc3, Amsterdamvarianten
D12.9=Slaviskt: 4.e3 Bf5 5.Bd3
D12.10=Slaviskt: 4.e3 Bf5 5.Bd3 Bxd3
D12.11=Slaviskt: 4.e3 Bf5 5.Nc3
D12.12=Slaviskt: 4.e3 Bf5 5.Nc3 e6
D12.13=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Be2
D12.14=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Bd3
D12.15=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Bd3 Bxd3
D12.16=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Bd3 Bxd3
D12.17=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Bd3 Bxd3 7.Qxd3 Nbd7
D12.18=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Nh4
D12.19=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Nh4 Bg4
D12.20=Slaviskt: 4.e3 Bf5 5.Nc3 e6 6.Nh4 Be4
D13.1=Slaviskt: Avbyte
D13.2=Slaviskt: Avbyte
D13.3=Slaviskt: Avbyte, 5.Nc3
D13.4=Slaviskt: Avbyte, 5.Nc3 Bf5
D13.5=Slaviskt: Avbyte, 5.Nc3 a6
D13.6=Slaviskt: Avbyte, 5.Nc3 a6 6.Ne5
D13.7=Slaviskt: Avbyte, 5.Nc3 a6 6.Bf4
D13.8=Slaviskt: Avbyte, 5.Nc3 e6
D13.9=Slaviskt: Avbyte, 5.Nc3 e6 6.Bf4
D13.10=Slaviskt: Avbyte, 5.Nc3 Nc6
D13.11=Slaviskt: Avbyte, 6.Bf4
D13.12=Slaviskt: Avbyte, 6.Bf4 a6
D13.13=Slaviskt: Avbyte, 6.Bf4 a6 7.e3
D13.14=Slaviskt: Avbyte, 6.Bf4 a6 7.e3 Bg4
D13.15=Slaviskt: Avbyte, 6.Bf4 a6 7.e3 Bg4 8.Be2
D13.16=Slaviskt: Avbyte, 6.Bf4 e6
D13.17=Slaviskt: Avbyte, 6.Bf4 e6 7.e3
D13.18=Slaviskt: Avbyte, 6.Bf4 e6 7.e3 Be7
D13.19=Slaviskt: Avbyte, 6.Bf4 e6 7.e3 Bd6
D13.20=Slaviskt: Avbyte, 6.Bf4 e6 7.e3 Bd6 8.Bxd6 Qxd6
D14.1=Slaviskt: Avbyte, 6.Bf4 Bf5
D14.2=Slaviskt: Avbyte, 6.Bf4 Bf5 7.e3
D14.3=Slaviskt: Avbyte, 6.Bf4 Bf5 7.e3 a6
D14.4=Slaviskt: Avbyte, 6.Bf4 Bf5 7.e3 e6
D14.5=Slaviskt: Avbyte, 8.Ne5
D14.6=Slaviskt: Avbyte, 8.Qb3
D14.7=Slaviskt: Avbyte, Trifunovicvarianten
D14.8=Slaviskt: Avbyte, 8.Bd3
D14.9=Slaviskt: Avbyte, 8.Bd3 Bxd3 9.Qxd3 Bd6
D14.10=Slaviskt: Avbyte, 8.Bd3 Bxd3 9.Qxd3 Bd6 10.Bxd6 Qxd6
D14.11=Slaviskt: Avbyte, 8.Bd3 Huvudvarianten
D14.12=Slaviskt: Avbyte, 8.Bd3 Huvudvarianten, 12.Rac1
D14.13=Slaviskt: Avbyte, 8.Bd3 Huvudvarianten, 12.Rfc1
D14.14=Slaviskt: Avbyte, 8.Bd3 Huvudvarianten, 12.Rfc1 Rfc8
D14.15=Slaviskt: Avbyte, 8.Bb5
D14.16=Slaviskt: Avbyte, 8.Bb5 Nd7
D14.17=Slaviskt: Avbyte, 8.Bb5 Nd7 9.Qa4
D15.1=Slaviskt: 4.Nc3
D15.2=Slaviskt: 4.Nc3 Bf5
D15.3=Slaviskt: 4.Nc3 Bf5 5.Qb3
D15.4=Slaviskt: S�chtingvarianten
D15.5=Slaviskt: Chameleonvarianten
D15.6=Slaviskt: Chameleon, 5.Bg5
D15.7=Slaviskt: Chameleon, 5.Ne5
D15.8=Slaviskt: Chameleon, 5.e3
D15.9=Slaviskt: Chameleon, 5.e3 b5
D15.10=Slaviskt: Chameleon, 5.e3 b5 6.b3
D15.11=Slaviskt: Chameleon, 5.c5
D15.12=Slaviskt: Chameleon, 5.c5 Nbd7
D15.13=Slaviskt: Chameleon, 5.a4
D15.14=Slaviskt: Chameleon, 5.a4 e6
D15.15=Slaviskt: Chameleon, 5.a4 e6 6.Bg5
D15.16=Slaviskt: Antagen
D15.17=Slaviskt: Antagen, 5.Ne5
D15.18=Slaviskt: Antagen, Alekhine
D15.19=Slaviskt: Antagen, Alekhine: 5...b5 6.a4 b4
D15.20=Slaviskt: Antagen, Alekhine: 5...b5 6.a4 b4 7.Nb1
D15.21=Slaviskt: Gellers (Tolush) gambit
D15.22=Slaviskt: Gellers gambit
D15.23=Slaviskt: Gellers gambit, Spasskyvarianten
D15.24=Slaviskt: Gellers gambit, 6.e5
D15.25=Slaviskt: Gellers gambit, 6.e5 Nd5 7.Ng5
D15.26=Slaviskt: Geller gambit, 6.e5 Nd5 7.a4
D15.27=Slaviskt: Gellers gambit, 6.e5 Nd5 7.a4 e6
D16.1=Slaviskt: Alapin
D16.2=Slaviskt: 5.a4 Nd5
D16.3=Slaviskt: Soultanbeieff-varianten
D16.4=Slaviskt: Mureyvarianten
D16.5=Slaviskt: Smyslovvarianten
D16.6=Slaviskt: Smyslov, 6.Ne5
D16.7=Slaviskt: Smyslov, 6.e3
D16.8=Slaviskt: Smyslov, 6.e3 Bg4
D16.9=Slaviskt: Smyslov, 6.e4
D16.10=Slaviskt: Smyslov, 6.e4 Bg4
D16.11=Slaviskt: Smyslov, 6.e4 Bg4 7.Bxc4 e6
D16.12=Slaviskt: Bronstein (Steiner)varianten
D16.13=Slaviskt: Bronstein, 6.Ne5
D16.14=Slaviskt: Bronstein, 6.Ne5 Bh5
D16.15=Slaviskt: Bronstein, 6.Ne5 Bh5 7.h3
D16.16=Slaviskt: Bronstein, 6.Ne5 Bh5 7.g3
D16.17=Slaviskt: Bronstein, 6.Ne5 Bh5 7.f3
D16.18=Slaviskt: Bronstein, 6.Ne5 Bh5 7.f3 Nfd7
D16.19=Slaviskt: Bronstein, 6.Ne5 Bh5 7.f3 Nfd7 8.Nxc4 e5 9.Ne4
D17.1=Slaviskt: Tjeckiskt f�rsvar
D17.2=Slaviskt: Tjeckiskt, 6.Nh4
D17.3=Slaviskt: Tjeckiskt, 6.Nh4 e6
D17.4=Slaviskt: Tjeckiskt, 6.Nh4 e6 7.Nxf5 exf5 8.e3
D17.5=Slaviskt: Tjeckiskt, 6.Nh4 Bc8
D17.6=Slaviskt: Tjeckiskt, 6.Nh4 Bc8 7.e3
D17.7=Slaviskt: Centrumvarianten
D17.8=Slaviskt: Centrum, 6.Ne5 Na6
D17.9=Slaviskt: Centrum, 6.Ne5 Na6 7.f3
D17.10=Slaviskt: Centrum, 6.Ne5 Nbd7
D17.11=Slaviskt: Centrum, Carlsbadvarianten
D17.12=Slaviskt: Centrum, Carlsbad, Huvudvarianten
D17.13=Slaviskt: Centrum, 6.Ne5 e6
D17.14=Slaviskt: Centrum, 6.Ne5 e6 7.f3
D17.15=Slaviskt: Centrum, H�bner (7...c5)
D17.16=Slaviskt: Centrum, 7.f3 Bb4
D17.17=Slaviskt: Centrum, 7.f3 Bb4 8.Bg5
D17.18=Slaviskt: Centrum, 7.f3 Bb4 8.Nxc4
D17.19=Slaviskt: Centrum, 7.f3 Bb4 8.e4
D17.20=Slaviskt: Centrum, Offra pj�s-varianten
D17.21=Slaviskt: Centrum, Huvudvarianten
D17.22=Slaviskt: Centrum, Huvudvarianten, 15.Nxc4
D17.23=Slaviskt: Centrum, Huvudvarianten, 15.Nxc4 O-O
D17.24=Slaviskt: Centrum, Huvudvarianten, 15.Nxc4 O-O-O
D18.1=Slaviskt: Holl�ndskta varianten
D18.2=Slaviskt: Holl�ndskt, Laskervarianten
D18.3=Slaviskt: Holl�ndskt, 6...e6
D18.4=Slaviskt: Holl�ndskt, 6...e6 7.Bxc4 Bb4
D18.5=Slaviskt: Holl�ndskt, 8.O-O
D18.6=Slaviskt: Holl�ndskt, 8...Nbd7
D18.7=Slaviskt: Holl�ndskt, 8...Nbd7 9.Nh4
D18.8=Slaviskt: Holl�ndskt, 8...Nbd7 9.Nh4 Bg6
D18.9=Slaviskt: Holl�ndskt, 8...Nbd7 9.Qb3
D18.10=Slaviskt: Holl�ndskt, 8...Nbd7 9.Qb3 a5
D18.11=Slaviskt: Holl�ndskt, 8...Nbd7 9.Qe2
D18.12=Slaviskt: Holl�ndskt, 8...Nbd7 9.Qe2 Bg6
D18.13=Slaviskt: Holl�ndskt, 8...Nbd7 9.Qe2 Bg6 10.e4
D18.14=Slaviskt: Holl�ndskt, 8...O-O
D18.15=Slaviskt: Holl�ndskt, 8...O-O 9.Qb3
D18.16=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4
D18.17=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Bg6
D18.18=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Bg4
D18.19=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Nbd7
D18.20=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Nbd7 10.Nxf5
D18.21=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Nbd7 10.Nxf5 exf5
D18.22=Slaviskt: Holl�ndskt, 8...O-O 9.Nh4 Nbd7 10.Nxf5 exf5 11.Qc2
D19.1=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2
D19.2=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg4
D19.3=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6
D19.4=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6 10.Rd1
D19.5=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6 10.Rd1 Nbd7
D19.6=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6 10.Ne5
D19.7=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6 10.Ne5 Nbd7, 12.Rd1
D19.8=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Bg6 10.Ne5 Nbd7, 12.Rd1
D19.9=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Ne4
D19.10=Slaviskt: Holl�ndskt, S�mischvarianten
D19.11=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7
D19.12=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4
D19.13=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg4
D19.14=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6
D19.15=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6 11.Bd3
D19.16=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6 11.Bd3 h6
D19.17=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6 11.Bd3 Re8
D19.18=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6 11.Bd3 Bh5
D19.19=Slaviskt: Holl�ndskt, 8...O-O 9.Qe2 Nbd7 10.e4 Bg6 11.Bd3 Bh5 12.e5
D20.1=Antagen damgambit
D20.2=Antagen damgambit: 3.Qa4+
D20.3=Antagen damgambit: 3.e3
D20.4=Antagen damgambit: 3.e3 c5
D20.5=Antagen damgambit: 3.e3 c5 4.Bxc4
D20.6=Antagen damgambit: 3.e3 c5 4.Bxc4
D20.7=Antagen damgambit: 3.e3 e6
D20.8=Antagen damgambit: 3.e3 e6
D20.9=Antagen damgambit: 3.e3 e5
D20.10=Antagen damgambit: 3.e3 e5
D20.11=Antagen damgambit: 3.e3 e5
D20.12=Antagen damgambit: 3.e3 e5
D20.13=Antagen damgambit: 3.e3 e5
D20.14=Antagen damgambit: 3.e3 Nf6
D20.15=Antagen damgambit: 3.Nc3
D20.16=Antagen damgambit: 3.Nc3 c5
D20.17=Antagen damgambit: 3.Nc3 e5
D20.18=Antagen damgambit: 3.Nc3 Nf6
D20.19=Antagen damgambit: 3.Nc3 e6
D20.20=Antagen damgambit: 3.Nc3 e6 4.e4
D20.21=Antagen damgambit: 3.Nc3 a6
D20.22=Antagen damgambit: 3.Nc3 a6 4.a4
D20.23=Antagen damgambit: 3.e4
D20.24=Antagen damgambit: 3.e4, Schwartz f�rsvar
D20.25=Antagen damgambit: 3.e4 Nc6
D20.26=Antagen damgambit: 3.e4 Nc6 4.Nf3
D20.27=Antagen damgambit: 3.e4 Nc6 4.Be3
D20.28=Antagen damgambit: 3.e4 Nf6
D20.29=Antagen damgambit: 3.e4 Nf6 4.Nc3
D20.30=Antagen damgambit: 3.e4 Nf6 4.e5
D20.31=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5
D20.32=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6
D20.33=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6 6.Bd3
D20.34=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6 6.Bd3
D20.35=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6 6.Bb3
D20.36=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6 6.Bb3
D20.37=Antagen damgambit: 3.e4 Nf6 4.e5 Nd5 5.Bxc4 Nb6 6.Bb3 Nc6 7.Ne2
D20.38=Antagen damgambit: 3.e4 c5
D20.39=Antagen damgambit: 3.e4 c5
D20.40=Antagen damgambit: 3.e4 c5 4.d5
D20.41=Antagen damgambit: Linaresvarianten
D20.42=Antagen damgambit: 3.e4 e5
D20.43=Antagen damgambit: 3.e4 e5 4.Nf3 Bb4+
D20.44=Antagen damgambit: 3.e4 e5 4.Nf3 exd4
D20.45=Antagen damgambit: 3.e4 e5 4.Nf3 exd4 5.Bxc4 Nc6
D21.1=Antagen damgambit: 3.Nf3
D21.2=Antagen damgambit: Ericsonvarianten
D21.3=Antagen damgambit: 3.Nf3 Nd7
D21.4=Antagen damgambit: 3.Nf3 Bg4
D21.5=Antagen damgambit: 3.Nf3 e6
D21.6=Antagen damgambit: 3.Nf3 e6 4.Qa4+
D21.7=Antagen damgambit: 3.Nf3 e6 4.e4
D21.8=Antagen damgambit: 3.Nf3 e6 4.e3
D21.9=Antagen damgambit: 3.Nf3 e6 4.e3 c5
D21.10=Antagen damgambit: 3.Nf3 c5
D21.11=Antagen damgambit: 3.Nf3 c5 4.Nc3
D21.12=Antagen damgambit: 3.Nf3 c5 4.e3
D21.13=Antagen damgambit: 3.Nf3 c5 4.e3 cxd4
D21.14=Antagen damgambit: 3.Nf3 c5 4.e3 cxd4 5.Bxc4
D21.15=Antagen damgambit: 3.Nf3 c5 4.d5
D21.16=Antagen damgambit: 3.Nf3 c5 4.d5 e6
D21.17=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.e4
D21.18=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.Nc3
D21.19=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.Nc3 exd5
D21.20=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.Nc3 exd5 6.Qxd5 Qxd5 7.Nxd5
D21.21=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.Nc3 exd5 6.Qxd5 Qxd5 7.Nxd5 Bd6
D21.22=Antagen damgambit: 3.Nf3 c5 4.d5 e6 5.Nc3 exd5 6.Qxd5 Qxd5 7.Nxd5 Bd6 8.Nd2
D21.23=Antagen damgambit: Seirawanvarianten
D21.24=Antagen damgambit: Alekhines f�rsvar
D21.25=Antagen damgambit: Alekhine, Borisenko-Furmanvarianten
D21.26=Antagen damgambit: Alekhine, 4.a4
D22.1=Antagen damgambit: Alekhine, 4.e3
D22.2=Antagen damgambit: Alekhine, Haberditzvarianten
D22.3=Antagen damgambit: Alekhine, 4.e3 e6
D22.4=Antagen damgambit: Alekhine, 4.e3 e6 5.Bxc4
D22.5=Antagen damgambit: Alekhine, 4.e3 e6 5.Bxc4 c5
D22.6=Antagen damgambit: Alekhine, 4.e3 e6 5.Bxc4 c5 6.Qe2
D22.7=Antagen damgambit: Alekhine, 4.e3 Bg4
D22.8=Antagen damgambit: Alekhine, 4.e3 Bg4 5.Bxc4 e6
D22.9=Antagen damgambit: Alekhine, Alatortsevvarianten
D22.10=Antagen damgambit: Alekhine, 4.e3 Bg4 5.Bxc4 e6 6.Qb3
D22.11=Antagen damgambit: Alekhine, 4.e3 Bg4 5.Bxc4 e6 6.Nc3
D22.12=Antagen damgambit: Alekhine, 4.e3 Bg4 5.Bxc4 e6 6.h3
D23.1=Antagen damgambit: 3.Nf3 Nf6
D23.2=Antagen damgambit: 3.Nf3 Nf6 4.g3
D23.3=Antagen damgambit: Mannheimvarianten
D23.4=Antagen damgambit: Mannheim, 4...Nc6
D23.5=Antagen damgambit: Mannheim, 4...Nc6
D23.6=Antagen damgambit: Mannheim, 4...Nbd7
D23.7=Antagen damgambit: Mannheim, 4...Nbd7 5.Nc3 e6
D23.8=Antagen damgambit: Mannheim, 4...Nbd7 5.Nc3 e6 6.e4
D23.9=Antagen damgambit: Mannheim, 4...c6
D23.10=Antagen damgambit: Mannheim, 4...c6 5.Qxc4
D23.11=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5
D23.12=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5 6.Nc3
D23.13=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5 6.g3
D23.14=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5 6.g3 e6
D23.15=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5 6.g3 e6 7.Bg2
D23.16=Antagen damgambit: Mannheim, 4...c6, 5.Qxc4 Bf5 6.g3 e6 7.Bg2 Nbd7
D23.17=Antagen damgambit: Mannheim, Huvudvarianten
D23.18=Antagen damgambit: Mannheim, Huvudvarianten, 9...O-O
D23.19=Antagen damgambit: Mannheim, Huvudvarianten, 10.Bg5
D23.20=Antagen damgambit: Mannheim, Huvudvarianten, 10.e3
D23.21=Antagen damgambit: Mannheim, Huvudvarianten, 10.e3 Ne4
D23.22=Antagen damgambit: Mannheim, Huvudvarianten, 10.e3 Ne4 11.Qe2
D24.1=Antagen damgambit: 4.Nc3
D24.2=Antagen damgambit: 4.Nc3 Nd5
D24.3=Antagen damgambit: 4.Nc3 e6
D24.4=Antagen damgambit: 4.Nc3 e6 5.Bg5
D24.5=Antagen damgambit: 4.Nc3 e6 5.e4
D24.6=Antagen damgambit: 4.Nc3 e6 5.e3
D24.7=Antagen damgambit: 4.Nc3 c5
D24.8=Antagen damgambit: 4.Nc3 c5 5.d5
D24.9=Antagen damgambit: 4.Nc3 c5 5.d5 e6 6.e4
D24.10=Antagen damgambit: 4.Nc3 c5 5.d5 e6 6.e4
D24.11=Antagen damgambit: 4.Nc3 c5 5.d5 e6 6.e4
D24.12=Antagen damgambit: 4.Nc3 c5 5.d5 e6 6.e4
D24.13=Antagen damgambit: 4.Nc3 a6
D24.14=Antagen damgambit: 4.Nc3 a6 5.a4
D24.15=Antagen damgambit: 4.Nc3 a6 5.a4 Nc6
D24.16=Antagen damgambit: 4.Nc3 a6 5.a4 Nc6 5.e4
D24.17=Antagen damgambit: Bogoljubow
D24.18=Antagen damgambit: Bogoljubow, 7.a4
D24.19=Antagen damgambit: Bogoljubow, 7.a4 e6
D24.20=Antagen damgambit: Bogoljubow, 7.a4 c6
D24.21=Antagen damgambit: Bogoljubow, 7.a4 Bb7
D24.22=Antagen damgambit: Bogoljubow, 7.a4 Nb4
D24.23=Antagen damgambit: Bogoljubow, 7.a4 Nxc3
D24.24=Antagen damgambit: Bogoljubow, 7.a4 Nxc3
D24.25=Antagen damgambit: Bogoljubow, 7.a4 Nxc3
D24.26=Antagen damgambit: Bogoljubow, 7.a4 Nxc3
D25.1=Antagen damgambit: 4.e3
D25.2=Antagen damgambit: 4.e3 c5
D25.3=Antagen damgambit: 4.e3 a6
D25.4=Antagen damgambit: Smyslovvarianten
D25.5=Antagen damgambit: Smyslov, 5.Bxc4 Bg7
D25.6=Antagen damgambit: Smyslov, 5.Bxc4 Bg7 6.O-O O-O
D25.7=Antagen damgambit: Flohrvarianten
D25.8=Antagen damgambit: Flohr, 5.Nc3
D25.9=Antagen damgambit: Flohr, 5.Nc3 c6
D25.10=Antagen damgambit: Janowski-Larsenvarianten
D25.11=Antagen damgambit: Janowski-Larsen, 5.h3
D25.12=Antagen damgambit: Janowski-Larsen, 5.Bxc4 e6
D25.13=Antagen damgambit: Janowski-Larsen, 6.Qb3
D25.14=Antagen damgambit: Janowski-Larsen, 6.O-O
D25.15=Antagen damgambit: Janowski-Larsen, 6.Nc3
D25.16=Antagen damgambit: Janowski-Larsen, 6.h3
D25.17=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3
D25.18=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 a6
D25.19=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 a6 8.g4
D25.20=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 Nbd7
D25.21=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 Nbd7 8.O-O
D25.22=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 Nbd7 8.O-O Bd6
D25.23=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 Nbd7 8.O-O Bd6 9.Be2
D25.24=Antagen damgambit: Janowski-Larsen, 6.h3 Bh5 7.Nc3 Nbd7 8.O-O Bd6 9.e4
D26.1=Antagen damgambit: 4.e3 e6
D26.2=Antagen damgambit: 4.e3 e6 5.Bxc4
D26.3=Antagen damgambit: 4.e3 e6 5.Bxc4 a6
D26.4=Antagen damgambit: 4.e3 e6 5.Bxc4 a6 6.O-O
D26.5=Antagen damgambit: 4.e3 e6 5.Bxc4 a6 6.O-O b5
D26.6=Antagen damgambit: Klassiska varianten
D26.7=Antagen damgambit: Klassisk, Tidigt dambyte
D26.8=Antagen damgambit: Klassisk, 6.Nc3
D26.9=Antagen damgambit: Klassisk, 6.Nc3 a6
D26.10=Antagen damgambit: Klassisk, Furmanvarianten
D26.11=Antagen damgambit: Klassisk, Furman, 6...cxd4
D26.12=Antagen damgambit: Klassisk, Furman, 6...a6
D26.13=Antagen damgambit: Klassisk, Furman, 6...a6 7.dxc5 Bxc5 8.O-O
D26.14=Antagen damgambit: Klassisk, Furman, 6...a6 7.dxc5 Bxc5 8.O-O Nc6
D26.15=Antagen damgambit: Klassisk, Furman, 6...a6 7.dxc5 Bxc5 8.O-O b5
D26.16=Antagen damgambit: Klassisk, 6.O-O
D26.17=Antagen damgambit: Klassisk, Steinitzvarianten
D26.18=Antagen damgambit: Klassisk, 6.O-O Nc6
D26.19=Antagen damgambit: Klassisk, 6.O-O Nc6 7.Nc3
D26.20=Antagen damgambit: Klassisk, 6.O-O Nc6 7.Qe2
D27.1=Antagen damgambit: Klassisk, 6...a6
D27.2=Antagen damgambit: Klassisk, 6...a6 7.a3
D27.3=Antagen damgambit: Klassisk, 6...a6 7.b3
D27.4=Antagen damgambit: Klassisk, 6...a6 7.Nc3
D27.5=Antagen damgambit: Klassisk, 6...a6 7.Bd3
D27.6=Antagen damgambit: Klassisk, 6...a6 7.Bd3 Nbd7
D27.7=Antagen damgambit: Klassisk, 6...a6 7.Bb3
D27.8=Antagen damgambit: Klassisk, 6...a6 7.Bb3 b5
D27.9=Antagen damgambit: Klassisk, 6...a6 7.Bb3 cxd4
D27.10=Antagen damgambit: Klassisk, 6...a6 7.Bb3 Nc6
D27.11=Antagen damgambit: Klassisk, 6...a6 7.Bb3 Nc6 8.Nc3
D27.12=Antagen damgambit: Klassisk, Gellervarianten
D27.13=Antagen damgambit: Klassisk, Spasskyvarianten
D27.14=Antagen damgambit: Klassisk, Spassky, 7...Qxd1
D27.15=Antagen damgambit: Klassisk, Spassky, 9.Nbd2
D27.16=Antagen damgambit: Klassisk, Spassky, 9.b3
D27.17=Antagen damgambit: Klassisk, Rubinsteinvarianten
D27.18=Antagen damgambit: Klassisk, Rubinstein, 7...Nc6
D27.19=Antagen damgambit: Klassisk, Rubinstein, 8.Nc3
D27.20=Antagen damgambit: Klassisk, Rubinstein, 8.Nc3 Be7
D27.21=Antagen damgambit: Klassisk, Rubinstein, 8.Nc3 Be7 9.Qe2
D27.22=Antagen damgambit: Klassisk, Rubinstein, 8.Qe2
D27.23=Antagen damgambit: Klassisk, Rubinstein, 8.Qe2 Qc7
D27.24=Antagen damgambit: Klassisk, Rubinstein, 8.Qe2 cxd4
D27.25=Antagen damgambit: Klassisk, Rubinstein, 8.Qe2 cxd4, 11.Nc3
D27.26=Antagen damgambit: Klassisk, Rubinstein, 8.Qe2 cxd4, 11.Nc3 Nd5
D28.1=Antagen damgambit: Klassisk, 7.Qe2
D28.2=Antagen damgambit: Klassisk, 7.Qe2 cxd4
D28.3=Antagen damgambit: Klassisk, 7.Qe2 Nc6
D28.4=Antagen damgambit: Klassisk, 7.Qe2 b5
D28.5=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bd3
D28.6=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bd3 cxd4
D28.7=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bd3 cxd4 9.exd4
D28.8=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3
D28.9=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6
D28.10=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6 9.Rd1
D28.11=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6 9.Rd1 c4
D28.12=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6 9.Nc3
D28.13=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6 9.Nc3 Bb7
D28.14=Antagen damgambit: Klassisk, 7.Qe2 b5 8.Bb3 Nc6 9.Nc3 Be7
D29.1=Antagen damgambit: Klassisk, 8...Bb7
D29.2=Antagen damgambit: Klassisk, 8...Bb7 9.Nc3
D29.3=Antagen damgambit: Klassisk, 8...Bb7 9.a4
D29.4=Antagen damgambit: Klassisk, 8...Bb7 9.a4 b4
D29.5=Antagen damgambit: Klassisk, 8...Bb7 9.a4 Nbd7
D29.6=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1
D29.7=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7
D29.8=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.e4
D29.9=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.a4
D29.10=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.a4 b4
D29.11=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.Nc3
D29.12=Antagen damgambit: Klassisk, Smyslovvarianten
D29.13=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.Nc3 Qc7
D29.14=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.Nc3 Qb8
D29.15=Antagen damgambit: Klassisk, 8...Bb7 9.Rd1 Nbd7 10.Nc3 Qb6
D30.1=Avb�jd damgambit)
D30.2=Avb�jd damgambit: 3.e3
D30.3=Diemer-Duhm gambit (DDG)
D30.4=Diemer-Duhm gambit (DDG) Antagen
D30.5=Diemer-Duhm gambit (DDG): 4...f5
D30.6=Diemer-Duhm gambit (DDG): Alapinvarianten
D30.7=Diemer-Duhm gambit (DDG): Duhmvarianten
D30.8=Diemer-Duhm gambit (DDG): 5.f3
D30.9=Diemer-Duhm gambit (DDG): Avbytesvarianten
D30.10=Diemer-Duhm gambit (DDG): Keres f�rsvar
D30.11=Diemer-Duhm gambit (DDG): Huvudvarianten
D30.12=Avb�jd damgambit: 3.g3
D30.13=Avb�jd damgambit: 3.cxd5
D30.14=Avb�jd damgambit: 3.cxd5
D30.15=Avb�jd damgambit: 3.cxd5
D30.16=Avb�jd damgambit: 3.Bf4
D30.17=Avb�jd damgambit: 3.Nf3
D30.18=Avb�jd damgambit: 3.Nf3 Nbd7 (Westphalia)
D30.19=Avb�jd damgambit: Tarrasch utan Nc3
D30.20=Avb�jd damgambit: Tarrasch utan Nc3: 4.e3
D30.21=Avb�jd damgambit: Tarrasch utan Nc3: 4.e3 Nf6
D30.22=Avb�jd damgambit: Tarrasch utan Nc3
D30.23=Avb�jd damgambit: Tarrasch utan Nc3
D30.24=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3
D30.25=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3
D30.26=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3
D30.27=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3 Nc6
D30.28=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3 Nc6 6.Bg2
D30.29=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3 Nc6 6.Bg2 Nf6
D30.30=Avb�jd damgambit: Tarrasch utan Nc3: 5.g3 Nc6 6.Bg2 Nf6 7.O-O
D30.31=Avb�jd damgambit: Tarrasch utan Nc3: Huvudvarianten
D30.32=Avb�jd damgambit: 3.Nf3 c6
D30.33=Avb�jd damgambit: 3.Nf3 c6 4.e3
D30.34=Avb�jd damgambit: 3.Nf3 c6 4.Nbd2
D30.35=Avb�jd damgambit: 3.Nf3 c6 4.Qc2
D30.36=Avb�jd damgambit: 3.Nf3 c6 4.Qc2 Nf6
D30.37=Avb�jd damgambit: 3.Nf3 c6 4.Qc2 Nf6 5.Bg5
D30.38=Avb�jd damgambit: 3.Nf3 c6 4.Qc2 Nf6 5.g3
D30.39=Avb�jd damgambit: 3.Nf3 Nf6
D30.40=Avb�jd damgambit: 3.Nf3 Nf6 4.e3
D30.41=Avb�jd damgambit: 3.Nf3 Nf6 4.e3 c6
D30.42=Avb�jd damgambit: 3.Nf3 Nf6 4.e3 c6 5.Nbd2
D30.43=Avb�jd damgambit: Spielmannvarianten
D30.44=Avb�jd damgambit: Stonewallformationen
D30.45=Avb�jd damgambit: 3.Nf3 Nf6 4.e3 c6 5.Nbd2 Nbd7
D30.46=Avb�jd damgambit: 3.Nf3 Nf6 4.e3 c6 5.Nbd2 Nbd7 6.Bd3
D30.47=Avb�jd damgambit: Semmeringvarianten
D30.48=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5
D30.49=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5 dxc4
D30.50=Avb�jd damgambit: Viennavarianten
D30.51=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5 Nbd7
D30.52=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5, Capablancavarianten
D30.53=Avb�jd damgambit: Capablanca-Duras varianten
D30.54=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5 Be7
D30.55=Avb�jd damgambit: 3.Nf3 Nf6 4.Bg5 Be7 5.e3
D31.1=Avb�jd damgambit: 3.Nc3
D31.2=Avb�jd damgambit: 3.Nc3 Nc6
D31.3=Avb�jd damgambit: Alapinvarianten
D31.4=Avb�jd damgambit: Janowskivarianten
D31.5=Avb�jd damgambit: 3.Nc3 Bb4
D31.6=Avb�jd damgambit: 3.Nc3 Bb4 4.a3
D31.7=Avb�jd damgambit: Alatortsevvarianten
D31.8=Avb�jd damgambit: Alatortsev, 4.Nf3
D31.9=Avb�jd damgambit: Alatortsev, 4.Bf4
D31.10=Avb�jd damgambit: Alatortsev, Avbyte
D31.11=Avb�jd damgambit: Alatortsev, Avbyte
D31.12=Avb�jd damgambit: Alatortsev, 5.Bf4
D31.13=Avb�jd damgambit: Alatortsev, 5.Bf4 c6
D31.14=Avb�jd damgambit: Alatortsev, 5.Bf4 c6 6.e3 Bf5
D31.15=Avb�jd damgambit: Alatortsev, 5.Bf4 c6 6.e3 Bf5 7.g4
D31.16=Semi-Slaviskt
D31.17=Semi-Slaviskt: 4.cxd5
D31.18=Semi-Slaviskt: 4.cxd5
D31.19=Semi-Slaviskt: 4.cxd5 exd5 5.Nf3
D31.20=Semi-Slaviskt: 4.cxd5 exd5 5.Nf3 Bf5
D31.21=Semi-Slaviskt: 4.cxd5 exd5 5.Bf4
D31.22=Semi-Slaviskt: 4.e3
D31.23=Semi-Slaviskt: 4.e3 Nf6
D31.24=Semi-Slaviskt: 4.Nf3
D31.25=Semi-Slaviskt: Noteboomvarianten
D31.26=Semi-Slaviskt: Noteboom, 5.a4
D31.27=Semi-Slaviskt: Noteboom, 5.a4 Bb4 6.e3 b5
D31.28=Semi-Slaviskt: Noteboom, Koomenvarianten
D31.29=Semi-Slaviskt: Noteboom, Jungevarianten
D31.30=Semi-Slaviskt: Noteboom, Abrahamsvarianten
D31.31=Semi-Slaviskt: Noteboom, Abrahams, Huvudvarianten
D31.32=Semi-Slaviskt: Noteboom, Abrahams, Huvudvarianten, 14.O-O O-O
D31.33=Semi-Slaviskt: Marshalls gambit
D31.34=Semi-Slaviskt: Marshalls gambit, 4...Bb4
D31.35=Semi-Slaviskt: Marshalls gambit, 4...dxe4
D31.36=Semi-Slaviskt: Marshalls gambit, Gunderams gambit
D31.37=Semi-Slaviskt: Marshalls gambit, 5.Nxe4
D31.38=Semi-Slaviskt: Marshalls gambit, 5.Nxe4 Nf6
D31.39=Semi-Slaviskt: Marshalls gambit, 5.Nxe4 Bb4+
D31.40=Semi-Slaviskt: Marshalls gambit, 5.Nxe4 Bb4+ 6.Nc3
D31.41=Semi-Slaviskt: Marshalls gambit, 5.Nxe4 Bb4+ 6.Bd2
D31.42=Semi-Slaviskt: Marshalls gambit, 8.Ne2
D31.43=Semi-Slaviskt: Marshalls gambit, 8.Be2
D31.44=Semi-Slaviskt: Marshalls gambit, 8.Be2 Na6
D32.1=Avb�jd damgambit Tarrasch
D32.2=Avb�jd damgambit Tarrasch: 4.e3
D32.3=Avb�jd damgambit Tarrasch: 4.Nf3
D32.4=Avb�jd damgambit Tarrasch: 4.Nf3 cxd4 5.Nxd4 e5
D32.5=Avb�jd damgambit Tarrasch: 4.cxd5
D32.6=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit
D32.7=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 5.Qxd4
D32.8=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 5.Qxd4 Nc6 6.Qd1 exd5 7.e3
D32.9=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 5.Qa4+
D32.10=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 7.Qxd5 Nc6
D32.11=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 7.Qxd5 Nc6 8.Bg5
D32.12=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, 7.Qxd5 Nc6 8.Nf3
D32.13=Avb�jd damgambit Tarrasch: von Hennig-Scharas gambit, Huvudvarianten (11.Be2 O-O-O)
D32.14=Avb�jd damgambit Tarrasch: 4.cxd5 exd5
D32.15=Avb�jd damgambit Tarrasch: 5.g3
D32.16=Avb�jd damgambit Tarrasch: 5.dxc5
D32.17=Avb�jd damgambit Tarrasch: 5.dxc5, Tarraschs gambit
D32.18=Avb�jd damgambit Tarrasch: Marshalls gambit
D32.19=Avb�jd damgambit Tarrasch: Marshalls gambit
D32.20=Avb�jd damgambit Tarrasch: Marshalls gambit, Modern 6.Bc4
D32.21=Avb�jd damgambit Tarrasch: Marshalls gambit, 6.d5
D32.22=Avb�jd damgambit Tarrasch: 5.Nf3
D32.23=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6
D32.24=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.Bf4
D32.25=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.Bf4 Nf6
D32.26=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.Bg5
D32.27=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.Bg5 Be7
D32.28=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3
D32.29=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6
D32.30=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Bb5
D32.31=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2
D32.32=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 Be7
D32.33=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 Be7 8.dxc5 Bxc5
D32.34=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 cxd4
D32.35=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 cxd4 8.Nxd4 Bd6
D32.36=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 cxd4 8.Nxd4 Bd6 9.O-O
D32.37=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 cxd4 8.Nxd4 Bd6 9.O-O O-O
D32.38=Avb�jd damgambit Tarrasch: 5.Nf3 Nc6 6.e3 Nf6 7.Be2 cxd4 8.Nxd4 Bd6 9.O-O O-O 10.b3
D33.1=Avb�jd damgambit Tarrasch: 6.g3 (Schlecter/Rubinstein)
D33.2=Avb�jd damgambit Tarrasch: 6.g3 cxd4
D33.3=Avb�jd damgambit Tarrasch: Svenska varianten
D33.4=Avb�jd damgambit Tarrasch: Svensk, Rey Ardid-varianten
D33.5=Avb�jd damgambit Tarrasch: Svensk, 7.Bg2
D33.6=Avb�jd damgambit Tarrasch: Svensk, 7.Bg2 Bb4 8.O-O Nge7
D33.7=Avb�jd damgambit Tarrasch: Svensk, 9.a3
D33.8=Avb�jd damgambit Tarrasch: Svensk, 9.Bd2
D33.9=Avb�jd damgambit Tarrasch: Svensk, 9.Ne5
D33.10=Avb�jd damgambit Tarrasch: Svensk, 9.e4
D33.11=Avb�jd damgambit Tarrasch: Svensk, 9.e4 dxe4
D33.12=Avb�jd damgambit Tarrasch: 6.g3 Nf6 (Prag)
D33.13=Avb�jd damgambit Tarrasch: 6.g3 Nf6 (Prag)
D33.14=Avb�jd damgambit Tarrasch: 7.Bg2 Be6
D33.15=Avb�jd damgambit Tarrasch: Wagnervarianten
D33.16=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4
D33.17=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4 8.Nxd4
D33.18=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4 8.Nxd4 Be7
D33.19=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4 8.Nxd4 Be7
D33.20=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4 8.Nxd4 Be7
D33.21=Avb�jd damgambit Tarrasch: 7.Bg2 cxd4 8.Nxd4 Be7 9.O-O O-O 10.Be3
D34.1=Avb�jd damgambit Tarrasch: 7.Bg2 Be7
D34.2=Avb�jd damgambit Tarrasch: 7.Bg2 Be7 8.O-O
D34.3=Avb�jd damgambit Tarrasch: 7.Bg2 Be7 8.O-O Be6
D34.4=Avb�jd damgambit Tarrasch: 8.O-O O-O (Huvudvarianten)
D34.5=Avb�jd damgambit Tarrasch: 9.b3
D34.6=Avb�jd damgambit Tarrasch: 9.b3 Ne4
D34.7=Avb�jd damgambit Tarrasch: 9.Bf4
D34.8=Avb�jd damgambit Tarrasch: 9.Be3
D34.9=Avb�jd damgambit Tarrasch: 9.dxc5
D34.10=Avb�jd damgambit Tarrasch: Tarraschs gambit
D34.11=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5
D34.12=Avb�jd damgambit Tarrasch: Retivarianten
D34.13=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5
D34.14=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5 Be6
D34.15=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5 Be6 11.Bxf6
D34.16=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5 d4
D34.17=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5 d4 11.Bxf6 Qxf6 12.Nd5
D34.18=Avb�jd damgambit Tarrasch: 9.dxc5 Bxc5 10.Bg5 d4 11.Bxf6: Huvudvarianten
D34.19=Avb�jd damgambit Tarrasch: 9.Bg5
D34.20=Avb�jd damgambit Tarrasch: 9.Bg5 Be6
D34.21=Avb�jd damgambit Tarrasch: Stoltzvarianten
D34.22=Avb�jd damgambit Tarrasch: Bogoljubowvarianten
D34.23=Avb�jd damgambit Tarrasch: 9.Bg5 c4
D34.24=Avb�jd damgambit Tarrasch: 9.Bg5 c4 10.Ne5 Be6 11.Nxc6
D34.25=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4
D34.26=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4
D34.27=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6
D34.28=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3
D34.29=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3 Re8
D34.30=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3 Re8 12.Qb3
D34.31=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3 Re8 12.Rc1
D34.32=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3 Re8 12.Rc1 Bf8
D34.33=Avb�jd damgambit Tarrasch: 9.Bg5 cxd4 10.Nxd4 h6 11.Be3 Re8 12.Rc1 Bf8 13.Nxc6
D35.1=Avb�jd damgambit: 3.Nc3 Nf6
D35.2=Avb�jd damgambit: 3.Nc3 Nf6 4.e3
D35.3=Avb�jd damgambit: Harrwitz attack
D35.4=Avb�jd damgambit: Katalansk utan Nf3
D35.5=Avb�jd damgambit: Avbyte
D35.6=Avb�jd damgambit: Avbyte, 4...Nxd5
D35.7=Avb�jd damgambit: Avbyte
D35.8=Avb�jd damgambit: Avbyte, S�mischvarianten
D35.9=Avb�jd damgambit: Avbyte, 5.Nf3
D35.10=Avb�jd damgambit: Avbyte, 5.Nf3 c6
D35.11=Avb�jd damgambit: Avbyte, 5.Nf3 c6 6.e3
D35.12=Avb�jd damgambit: Avbyte, 5.Nf3 Nbd7
D35.13=Avb�jd damgambit: Avbyte, 5.Nf3 Nbd7 6.e3
D35.14=Avb�jd damgambit: Avbyte, 5.Nf3 Nbd7 6.e3 c6
D35.15=Avb�jd damgambit: Avbyte, 5.Nf3 Nbd7 6.Bf4
D35.16=Avb�jd damgambit: Avbyte, 5.Nf3 Be7
D35.17=Avb�jd damgambit: Avbyte, 5.Nf3 Be7 6.Bf4
D35.18=Avb�jd damgambit: Avbyte, 5.Nf3 Be7 6.Bf4 c6
D35.19=Avb�jd damgambit: Avbyte, 5.Nf3 Be7 6.Bf4 c6 7.Qc2
D35.20=Avb�jd damgambit: Avbyte, 5.Nf3 Be7 6.Bf4 c6 7.Qc2 Nbd7
D35.21=Avb�jd damgambit: Avbyte, 5.Bg5
D35.22=Avb�jd damgambit: Avbyte, 5.Bg5 Nbd7
D35.23=Avb�jd damgambit: Avbyte, 5.Bg5 Nbd7 6.Nf3
D35.24=Avb�jd damgambit: Avbyte, 5.Bg5 Nbd7 6.e3
D35.25=Avb�jd damgambit: Avbyte, 5.Bg5 Be7
D35.26=Avb�jd damgambit: Avbyte, 5.Bg5 Be7 6.Nf3
D35.27=Avb�jd damgambit: Avbyte, 5.Bg5 Be7 6.e3
D35.28=Avb�jd damgambit: Avbyte, 5.Bg5 Be7 6.e3 h6
D35.29=Avb�jd damgambit: Avbyte, 5.Bg5 Be7 6.e3 Nbd7
D35.30=Avb�jd damgambit: Avbyte, 5.Bg5 Be7 6.e3 O-O
D35.31=Avb�jd damgambit: Avbyte, 5.Bg5 c6
D35.32=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.Nf3
D35.33=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3
D35.34=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Nbd7
D35.35=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7
D35.36=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Nf3
D35.37=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Nf3 Bf5
D35.38=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Nf3 Bf5 8.Bd3
D35.39=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3
D35.40=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 Ne4
D35.41=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 Nbd7
D35.42=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 Nbd7 8.Nge2
D35.43=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 Nbd7 8.Nf3
D35.44=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 O-O
D35.45=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 O-O 8.Nf3
D35.46=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.e3 Be7 7.Bd3 O-O 8.Nge2
D36.1=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.Qc2
D36.2=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.Qc2 g6
D36.3=Avb�jd damgambit: Avbyte, 5.Bg5 c6 6.Qc2 Na6
D36.4=Avb�jd damgambit: Avbyte, 6.Qc2 Be7
D36.5=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.Nf3
D36.6=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.Nf3 Nbd7
D36.7=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.Nf3 O-O
D36.8=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.Nf3 g6
D36.9=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.Nf3 g6 8.e3
D36.10=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3
D36.11=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 O-O
D36.12=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 O-O 8.Bd3
D36.13=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 h6
D36.14=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 h6
D36.15=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 h6
D36.16=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 Nbd7
D36.17=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 Nbd7 8.Nf3
D36.18=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 Nbd7 8.Bd3
D36.19=Avb�jd damgambit: Avbyte, 6.Qc2 Be7 7.e3 Nbd7 8.Bd3 Nf8
D36.20=Avb�jd damgambit: Avbyte, Huvudvarianten
D36.21=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2
D36.22=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 h6
D36.23=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 h6 10.Bh4
D36.24=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 Re8
D36.25=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 Re8 10.O-O
D36.26=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 Re8 10.O-O Nf8
D36.27=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nge2 Re8 10.O-O Nf8 11.f3
D36.28=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3
D36.29=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 h6
D36.30=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 h6 10.Bh4
D36.31=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8
D36.32=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.h3
D36.33=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.h3 Nf8
D36.34=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.h3 Nf8 11.Bf4
D36.35=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O-O
D36.36=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O-O h6
D36.37=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O-O Nf8
D36.38=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O-O Nf8 11.h3
D36.39=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O
D36.40=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O h6
D36.41=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O h6
D36.42=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O h6
D36.43=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8
D36.44=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8 11.Rae1
D36.45=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8 11.h3
D36.46=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8 11.h3 g6
D36.47=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8 11.Rab1
D36.48=Avb�jd damgambit: Avbyte, Huvudvarianten, 9.Nf3 Re8 10.O-O Nf8 11.Rab1 a5
D37.1=Avb�jd damgambit: 4.Nf3
D37.2=Avb�jd damgambit: Westphalia utan Bg5
D37.3=Avb�jd damgambit: Westphalia: 4.Nf3 Nbd7 5.Bf4
D37.4=Avb�jd damgambit: 4.Nf3 Be7
D37.5=Avb�jd damgambit: 4.Nf3 Be7 5.cxd5 Nxd5
D37.6=Avb�jd damgambit: 4.Nf3 Be7 5.e3
D37.7=Avb�jd damgambit: 4.Nf3 Be7 5.e3 O-O
D37.8=Avb�jd damgambit: 4.Nf3 Be7 5.e3 O-O 6.b3
D37.9=Avb�jd damgambit: 4.Nf3 Be7 5.e3 O-O 6.Bd3
D37.10=Avb�jd damgambit: Klassiska varianten
D37.11=Avb�jd damgambit: Klassisk, 5...O-O
D37.12=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 Nbd7
D37.13=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 b6
D37.14=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c6
D37.15=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5
D37.16=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5
D37.17=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5
D37.18=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.a3
D37.19=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.cxd5
D37.20=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.Qc2
D37.21=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.Qc2 Nc6 9.a3
D37.22=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.Qc2 Nc6 9.a3 Qa5
D37.23=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.Qc2 Nc6 9.a3 Qa5 10.Rd1
D37.24=Avb�jd damgambit: Klassisk, 5...O-O 6.e3 c5 7.dxc5 Bxc5 8.Qc2 Nc6 9.a3 Qa5 10.O-O-O
D38.1=Avb�jd damgambit: Ragozin
D38.2=Avb�jd damgambit: Ragozin, 5.Qa4+
D38.3=Avb�jd damgambit: Ragozin, 5.Qa4+ Nc6 6.cxd5
D38.4=Avb�jd damgambit: Ragozin, 5.Qa4+ Nc6 6.cxd5 exd5 7.Bg5
D38.5=Avb�jd damgambit: Ragozin, 5.cxd5
D38.6=Avb�jd damgambit: Ragozin, 5.cxd5 exd5 6.Bg5
D38.7=Avb�jd damgambit: Ragozin, 5.cxd5 exd5 6.Bg5 h6
D38.8=Avb�jd damgambit: Ragozin, 5.cxd5 exd5 6.Bg5 h6
D38.9=Avb�jd damgambit: Ragozin, 5.Bg5
D38.10=Avb�jd damgambit: Ragozin, Westphalia-varianten
D38.11=Avb�jd damgambit: Ragozin, Westphalia, 7.Qc2
D38.12=Avb�jd damgambit: Ragozin, Westphalia, 7.e3
D38.13=Avb�jd damgambit: Ragozin, 5.Bg5 h6
D38.14=Avb�jd damgambit: Ragozin, 5.Bg5 h6 6.Bxf6 Qxf6
D38.15=Avb�jd damgambit: Ragozin, 5.Bg5 h6 6.Bxf6 Qxf6 7.cxd5
D38.16=Avb�jd damgambit: Ragozin, 5.Bg5 h6 6.Bxf6 Qxf6 7.cxd5
D38.17=Avb�jd damgambit: Ragozin, 5.Bg5 h6 6.Bxf6 Qxf6 7.e3
D38.18=Avb�jd damgambit: Ragozin, 5.Bg5 h6 6.Bxf6 Qxf6 7.e3 O-O 8.Rc1
D39.1=Avb�jd damgambit: Ragozin, Vienna-varianten
D39.2=Avb�jd damgambit: Ragozin, Vienna, 6.Qa4+
D39.3=Avb�jd damgambit: Ragozin, Vienna, 6.e4
D39.4=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5
D39.10=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.e5
D39.11=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.e5 cxd4
D39.12=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.e5 cxd4 8.Qa4+ Nc6 9.O-O-O
D39.5=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.Bxc4
D39.6=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.Bxc4
D39.7=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.Bxc4
D39.8=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.Bxc4, 8...Qa5
D39.9=Avb�jd damgambit: Ragozin, Vienna, 6.e4 c5 7.Bxc4, 8...Bxc3+
D40.1=Avb�jd damgambit: Semi-Tarrasch
D40.2=Avb�jd damgambit: Semi-Tarrasch, 5.e3
D40.3=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Be7
D40.4=Avb�jd damgambit: Semi-Tarrasch, 5.e3 cxd4
D40.5=Avb�jd damgambit: Semi-Tarrasch, 5.e3 a6
D40.6=Avb�jd damgambit: Semi-Tarrasch, 5.e3 a6 6.cxd5
D40.7=Avb�jd damgambit: Semi-Tarrasch, 5.e3 a6 6.cxd5 exd5
D40.8=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6
D40.9=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.Bd3
D40.10=Avb�jd damgambit: Semi-Tarrasch, Symmetriska varianten
D40.11=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3
D40.12=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 Ne4
D40.13=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 dxc4
D40.14=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 cxd4
D40.15=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 cxd4 7.exd4 Be7
D40.16=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 cxd4 7.exd4 Be7 8.c5
D40.17=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 cxd4 7.exd4 Be7 8.Bd3
D40.18=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 a6
D40.19=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 a6 7.b3
D40.20=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 a6 7.dxc5
D40.21=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 a6 7.dxc5 Bxc5
D40.22=Avb�jd damgambit: Semi-Tarrasch, 5.e3 Nc6 6.a3 a6 7.dxc5 Bxc5 8.b4 Ba7
D41.1=Avb�jd damgambit: Semi-Tarrasch, 5.cxd5
D41.2=Avb�jd damgambit: Semi-Tarrasch, Keres motattack
D41.3=Avb�jd damgambit: Semi-Tarrasch, 5.cxd5 Nxd5
D41.4=Avb�jd damgambit: Semi-Tarrasch, 6.g3
D41.5=Avb�jd damgambit: Semi-Tarrasch, 6.g3 Nc6
D41.6=Avb�jd damgambit: Semi-Tarrasch, 6.g3 Nc6 7.Bg2 Be7
D41.7=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten
D41.8=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.e4
D41.9=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.e4 Nb6
D41.10=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.e4 Ndb4
D41.11=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.Nxd5
D41.12=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.Nxd5 exd5 10.dxc5 Bxc5
D41.13=Avb�jd damgambit: Semi-Tarrasch, 6.g3, Huvudvarianten, 9.Nxd5 exd5 10.dxc5 Bxc5 11.Bg5
D41.14=Avb�jd damgambit: Semi-Tarrasch, 6.e4
D41.15=Avb�jd damgambit: Semi-Tarrasch, 6.e4 Nxc3
D41.16=Avb�jd damgambit: Semi-Tarrasch, 6.e4, 8.cxd4
D41.17=Avb�jd damgambit: Semi-Tarrasch, 6.e4, 8.cxd4 Nc6
D41.18=Avb�jd damgambit: Semi-Tarrasch, 6.e4, 8.cxd4 Bb4+
D41.19=Avb�jd damgambit: Semi-Tarrasch, 6.e4, San Sebastian-varianten
D41.20=Avb�jd damgambit: Semi-Tarrasch, 6.e4, Kmochvarianten
D41.21=Avb�jd damgambit: Semi-Tarrasch, 6.e4, Huvudvarianten
D41.22=Avb�jd damgambit: Semi-Tarrasch, 6.e4, Huvudvarianten
D41.23=Avb�jd damgambit: Semi-Tarrasch, 6.e4, Huvudvarianten, 12...b6
D41.24=Avb�jd damgambit: Semi-Tarrasch, 6.e4, Huvudvarianten, 12...b6
D41.25=Avb�jd damgambit: Semi-Tarrasch, 6.e3
D41.26=Avb�jd damgambit: Semi-Tarrasch, 6.e3 cxd4
D41.27=Avb�jd damgambit: Semi-Tarrasch, 6.e3 cxd4 7.exd4
D41.28=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6
D41.29=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bc4
D41.30=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bc4
D41.31=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bc4
D41.32=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bc4
D41.33=Avb�jd damgambit: Semi-Tarrasch, 7.Bc4 Huvudvarianten
D41.34=Avb�jd damgambit: Semi-Tarrasch, 7.Bc4 Huvudvarianten
D41.35=Avb�jd damgambit: Semi-Tarrasch, 7.Bc4 Huvudvarianten, 13.Qc2
D41.36=Avb�jd damgambit: Semi-Tarrasch, 7.Bc4 Huvudvarianten, 13.h4
D42.1=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bd3
D42.2=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bd3 Be7
D42.3=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bd3 Be7 8.O-O O-O
D42.4=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bd3 cxd4
D42.5=Avb�jd damgambit: Semi-Tarrasch, 6.e3 Nc6 7.Bd3 cxd4
D42.6=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten
D42.7=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 9.O-O O-O
D42.8=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.a3
D42.9=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.a3 Nf6
D42.10=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.a3 Bf6
D42.11=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1
D42.12=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Ncb4
D42.13=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6
D42.14=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.Bg5
D42.15=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.a3
D42.16=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.a3 b6
D42.17=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.a3 b6 12.Be3
D42.18=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.a3 b6 12.Bg5
D42.19=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Nf6 11.a3 b6 12.Bc2
D42.20=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Bf6
D42.21=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Bf6 11.Be4
D42.22=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Bf6 11.Be4 Nce7
D42.23=Avb�jd damgambit: Semi-Tarrasch, 7.Bd3 Huvudvarianten, 10.Re1 Bf6 11.Be4 Nce7 12.Ne5
D43.1=Semi-Slaviskt
D43.2=Semi-Slaviskt: 5.g3
D43.3=Semi-Slaviskt: 5.Qd3
D43.4=Semi-Slaviskt: 5.Qb3
D43.5=Semi-Slaviskt: 5.Qb3 dxc4
D43.6=Semi-Slaviskt: Botvinnik (Anti-Meran)
D43.7=Semi-Slaviskt: Botvinnik, 5...Be7
D43.8=Semi-Slaviskt: Botvinnik, 5...Be7 6.e3
D43.9=Semi-Slaviskt: Botvinnik, 5...Be7 6.e3 O-O
D43.10=Semi-Slaviskt: Botvinnik, 5...Be7 6.e3 Nbd7
D43.11=Semi-Slaviskt: Botvinnik, 5...Be7 6.e3 Nbd7 7.Bd3
D43.12=Semi-Slaviskt: Moskvavarianten
D43.13=Semi-Slaviskt: Moskva, 6.Bh4 gambit
D43.14=Semi-Slaviskt: Moskva, 6.Bh4 Be7
D43.15=Semi-Slaviskt: Moskva, 6.Bh4 Be7 7.e3 O-O
D43.16=Semi-Slaviskt: Antagen Moskva, 6.Bh4 gambit
D43.17=Semi-Slaviskt: Moskva, 6.Bh4 gambit, 7.e4
D43.18=Semi-Slaviskt: Moskva, 6.Bh4 gambit, Huvudvarianten
D43.19=Semi-Slaviskt: Moskva, 6.Bh4 gambit, Huvudvarianten, 9...Bb7
D43.20=Semi-Slaviskt: Moskva, 6.Bxf6
D43.21=Semi-Slaviskt: Moskva, 7.g3
D43.22=Semi-Slaviskt: Moskva, Hastingsvarianten
D43.23=Semi-Slaviskt: Moskva, 7.Qc2
D43.24=Semi-Slaviskt: Moskva, 7.e3
D43.25=Semi-Slaviskt: Moskva, 7.e3 Nd7
D43.26=Semi-Slaviskt: Moskva, 7.e3 Nd7 8.Bd3
D43.27=Semi-Slaviskt: Moskva, 7.e3 Nd7 8.Bd3 dxc4
D43.28=Semi-Slaviskt: Moskva, Huvudvarianten
D43.29=Semi-Slaviskt: Moskva, Huvudvarianten
D43.30=Semi-Slaviskt: Moskva, Huvudvarianten
D43.31=Semi-Slaviskt: Moskva, Huvudvarianten, 11.b4
D43.32=Semi-Slaviskt: Moskva, Huvudvarianten, 11.Rc1
D44.1=Semi-Slaviskt: Antagen Botvinnik
D44.2=Semi-Slaviskt: Botvinnik, 6.a4
D44.3=Semi-Slaviskt: Botvinnik, 6.e4
D44.4=Semi-Slaviskt: Botvinnik, 6.e4
D44.5=Semi-Slaviskt: Botvinnik, 7.a4
D44.6=Semi-Slaviskt: Botvinnik, 7.e5
D44.7=Semi-Slaviskt: Botvinnik, 9.exf6
D44.8=Semi-Slaviskt: Botvinnik, Ekstr�ms-varianten
D44.9=Semi-Slaviskt: Botvinnik, 9.Nxg5
D44.10=Semi-Slaviskt: Botvinnik, Alatortse-varianten
D44.11=Semi-Slaviskt: Botvinnik, 9.Nxg5
D44.12=Semi-Slaviskt: Botvinnik, Lilienthal-varianten
D44.13=Semi-Slaviskt: Botvinnik, Lilienthal, 11...Qa5
D44.14=Semi-Slaviskt: Botvinnik, Lilienthal, 11...Bb7
D44.15=Semi-Slaviskt: Botvinnik, Szabovarianten
D44.16=Semi-Slaviskt: Botvinnik, Huvudvarianten
D44.17=Semi-Slaviskt: Botvinnik, Huvudvarianten, 12.g3
D44.18=Semi-Slaviskt: Botvinnik, Huvudvarianten, 12.g3 c5
D44.19=Semi-Slaviskt: Botvinnik, Huvudvarianten, 12.g3 c5 13.d5 Qb6
D45.1=Semi-Slaviskt: 5.e3
D45.2=Semi-Slaviskt: 5.e3 Bd6
D45.3=Semi-Slaviskt: 5.e3 Be7
D45.4=Semi-Slaviskt: 5.e3 Ne4
D45.5=Semi-Slaviskt: Stonewallf�rsvar
D45.6=Semi-Slaviskt: Accelererad Meran (Alekhinevarianten)
D45.7=Semi-Slaviskt: 5.e3 Nbd7
D45.8=Semi-Slaviskt: Rubinsteins system
D45.9=Semi-Slaviskt: 6.a3
D45.10=Semi-Slaviskt: 6.Qc2
D45.11=Semi-Slaviskt: 6.Qc2 b6
D45.12=Semi-Slaviskt: 6.Qc2 Be7
D45.13=Semi-Slaviskt: 6.Qc2 Bd6
D45.14=Semi-Slaviskt: 6.Qc2 Bd6 7.e4
D45.15=Semi-Slaviskt: 6.Qc2 Bd6 7.g4
D45.16=Semi-Slaviskt: 6.Qc2 Bd6 7.g4 h6
D45.17=Semi-Slaviskt: 6.Qc2 Bd6 7.g4 dxc4
D45.18=Semi-Slaviskt: 6.Qc2 Bd6 7.g4 Bb4
D45.19=Semi-Slaviskt: 6.Qc2 Bd6 7.g4 Nxg4
D45.20=Semi-Slaviskt: 6.Qc2 Bd6 7.b3
D45.21=Semi-Slaviskt: 6.Qc2 Bd6 7.b3 O-O
D45.22=Semi-Slaviskt: 6.Qc2 Bd6 7.b3 O-O 8.Bb2
D45.23=Semi-Slaviskt: 6.Qc2 Bd6 7.b3 O-O 8.Be2
D45.24=Semi-Slaviskt: 6.Qc2 Bd6 7.b3 O-O 8.Be2 b6
D45.25=Semi-Slaviskt: 6.Qc2 Bd6 7.b3 O-O 8.Be2 Re8
D45.26=Semi-Slaviskt: 6.Qc2 Bd6 7.Bd2
D45.27=Semi-Slaviskt: 6.Qc2 Bd6 7.Be2
D45.28=Semi-Slaviskt: 6.Qc2 Bd6 7.Be2 O-O 8.O-O
D45.29=Semi-Slaviskt: 6.Qc2 Bd6 7.Be2 O-O 8.O-O e5
D45.30=Semi-Slaviskt: 6.Qc2 Bd6 7.Be2 O-O 8.O-O Qe7
D45.31=Semi-Slaviskt: 6.Qc2 Bd6 7.Be2 O-O 8.O-O Re8
D46.1=Semi-Slaviskt: 6.Bd3
D46.2=Semi-Slaviskt: 6.Bd3 a6
D46.3=Semi-Slaviskt: Romihvarianten
D46.4=Semi-Slaviskt: Romih, 7.O-O
D46.5=Semi-Slaviskt: Romih, 7.O-O O-O
D46.6=Semi-Slaviskt: Bogoljubowvarianten
D46.7=Semi-Slaviskt: Bogoljubow, 7.O-O
D46.8=Semi-Slaviskt: Bogoljubow, 7.O-O O-O
D46.9=Semi-Slaviskt: Bogoljubow, 7.O-O O-O 8.b3
D46.10=Semi-Slaviskt: Chigorins f�rsvar
D46.11=Semi-Slaviskt: Chigorin, 7.e4
D46.12=Semi-Slaviskt: Chigorin, 7.e4 dxe4 8.Nxe4
D46.13=Semi-Slaviskt: Chigorin, 7.Qc2
D46.14=Semi-Slaviskt: Chigorin, 7.Qc2 dxc4
D46.15=Semi-Slaviskt: Chigorin, 7.Qc2 dxc4
D46.16=Semi-Slaviskt: Chigorin, 7.Qc2 O-O
D46.17=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten
D46.18=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...e5
D46.19=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...Qe7
D46.20=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...Qe7 10.Bd2
D46.21=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...Qe7 10.a3
D46.22=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...Qe7 10.h3
D46.23=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...a6
D46.24=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...a6 10.Rd1
D46.25=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...a6 10.Rd1 b5
D46.26=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...b5
D46.27=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...b5 10.Be2
D46.28=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...b5 10.Be2 Bb7
D46.29=Semi-Slaviskt: Chigorin, 7.Qc2 Huvudvarianten, 9...b5 10.Be2 Bb7 11.Rd1
D46.30=Semi-Slaviskt: Chigorin, 7.O-O
D46.31=Semi-Slaviskt: Chigorin, 7.O-O O-O
D46.32=Semi-Slaviskt: Chigorin, 7.O-O O-O 8.e4
D46.33=Semi-Slaviskt: Chigorin, 7.O-O O-O 8.e4 dxc4
D46.34=Semi-Slaviskt: Chigorin, 7.O-O O-O 8.e4 dxc4 9.Bxc4
D46.35=Semi-Slaviskt: Chigorin, 7.O-O O-O 8.e4 dxc4 9.Bxc4 e5
D46.36=Semi-Slaviskt: Chigorin, Huvudvarianten
D46.37=Semi-Slaviskt: Chigorin, Huvudvarianten
D46.38=Semi-Slaviskt: Chigorin, Huvudvarianten
D46.39=Semi-Slaviskt: Chigorin, Huvudvarianten, 10...h6
D46.40=Semi-Slaviskt: Chigorin, Huvudvarianten, 10...h6 11.Bc2
D46.41=Semi-Slaviskt: Chigorin, Huvudvarianten, 10...h6 11.Bc2 e5
D47.1=Semi-Slaviskt: Meranvarianten
D47.2=Semi-Slaviskt: Meranvarianten
D47.3=Semi-Slaviskt: Meran, 7...b5
D47.4=Semi-Slaviskt: Meran, Freymannvarianten
D47.5=Semi-Slaviskt: Meran, Freymann, 8...b4
D47.6=Semi-Slaviskt: Meran, Capablancavarianten
D47.7=Semi-Slaviskt: Meran, Capablanca, 8...b4
D47.8=Semi-Slaviskt: Meran, Capablanca, 8...a6
D47.9=Semi-Slaviskt: Meran, Capablanca, 8...Bb7
D47.10=Semi-Slaviskt: Meran, Capablanca, 8...Bb7 9.O-O
D47.11=Semi-Slaviskt: Meran, Capablanca, 8...Bb7 9.O-O a6
D47.12=Semi-Slaviskt: Meran, 8.Bd3
D47.13=Semi-Slaviskt: Meran, 8.Bd3 Bd6
D47.14=Semi-Slaviskt: Meran, Lundinvarianten
D47.15=Semi-Slaviskt: Meran, Lundin, 9.Na4
D47.16=Semi-Slaviskt: Meran, Lundin, 9.Ne4
D47.17=Semi-Slaviskt: Meran, Lundin, 9.Ne4 Nxe4
D47.18=Semi-Slaviskt: Meran, Lundin, 9.Ne4 Be7
D47.19=Semi-Slaviskt: Meran, Lundin, 9.Ne4 Be7 10.O-O
D47.20=Semi-Slaviskt: Meran, Wadevarianten
D47.21=Semi-Slaviskt: Meran, Wade, 9.a3
D47.22=Semi-Slaviskt: Meran, Wade, 9.O-O
D47.23=Semi-Slaviskt: Meran, Wade, 9.O-O b4
D47.24=Semi-Slaviskt: Meran, Wade, 9.O-O b4 10.Ne4
D47.25=Semi-Slaviskt: Meran, Wade, 9.O-O b4 10.Ne4 Be7
D47.26=Semi-Slaviskt: Meran, Wade, 9.O-O b4 10.Ne4 Be7 11.Nxf6+
D47.27=Semi-Slaviskt: Meran, Wade, 9.O-O b4 10.Ne4 Be7 11.Nxf6+ Nxf6
D47.28=Semi-Slaviskt: Meran, Wade, 9.O-O b4 10.Ne4 Be7 11.Nxf6+ Nxf6 12.e4
D47.29=Semi-Slaviskt: Meran, Wade, 9.e4
D47.30=Semi-Slaviskt: Meran, Wade, Huvudvarianten
D47.31=Semi-Slaviskt: Meran, Wade, Huvudvarianten, 12.Nxc5
D47.32=Semi-Slaviskt: Meran, Wade, Huvudvarianten, 12.O-O
D48.1=Semi-Slaviskt: Meran, 8...a6
D48.2=Semi-Slaviskt: Meran, 8...a6 9.a4
D48.3=Semi-Slaviskt: Meran, 8...a6 9.O-O
D48.4=Semi-Slaviskt: Meran, 8...a6 9.O-O c5
D48.5=Semi-Slaviskt: Meran, 8...a6 9.O-O c5 10.Qe2
D48.6=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7
D48.7=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7 10.e4
D48.8=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7 10.e4 c5 11.d5
D48.9=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7 10.e4 c5 11.d5 Qc7
D48.10=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7 10.e4 c5 11.d5 Qc7 12.dxe6
D48.11=Semi-Slaviskt: Meran, 8...a6 9.O-O Bb7 10.e4 c5 11.d5 Qc7 12.dxe6 fxe6
D48.12=Semi-Slaviskt: Meran, 8...a6 9.e4
D48.13=Semi-Slaviskt: Meran, 8...a6 9.e4 Bb7
D48.14=Semi-Slaviskt: Meran, Pircvarianten
D48.15=Semi-Slaviskt: Meran, 8...a6 9.e4 c5
D48.16=Semi-Slaviskt: Meran, Reynoldvarianten
D48.17=Semi-Slaviskt: Meran, Reynolds, 10...e5
D48.18=Semi-Slaviskt: Meran, Reynolds, 10...Qc7
D48.19=Semi-Slaviskt: Meran, Reynolds, 10...c4
D48.20=Semi-Slaviskt: Meran, Reynolds, 10...c4 11.dxe6 fxe6
D48.21=Semi-Slaviskt: Meran, Reynolds, 10...c4 11.dxe6 fxe6 12.Bc2
D48.22=Semi-Slaviskt: Meran, Reynolds, 10...c4 11.dxe6 fxe6 12.Bc2 Qc7
D48.23=Semi-Slaviskt: Meran, Reynolds, 10...c4 11.dxe6 fxe6 12.Bc2 Qc7 13.O-O
D48.24=Semi-Slaviskt: Meran, Gamla Huvudvarianten
D48.25=Semi-Slaviskt: Meran, Rabinovichvarianten
D48.26=Semi-Slaviskt: Meran, Gamla Huvudvarianten, 10...cxd4
D49.1=Semi-Slaviskt: Meran, Blumenfeldvarianten
D49.2=Semi-Slaviskt: Meran, Gamla Huvudvarianten, Gligoricvarianten
D49.3=Semi-Slaviskt: Meran, Gamla Huvudvarianten, Gligoric, 12.Qa4
D49.4=Semi-Slaviskt: Meran, Trifunovicvarianten
D49.5=Semi-Slaviskt: Meran, Sozinvarianten
D49.6=Semi-Slaviskt: Meran, Sozin, Rellstabattacken
D49.7=Semi-Slaviskt: Meran, Sozin, St�hlbergattacken
D49.8=Semi-Slaviskt: Meran, Sozin, St�hlbergattacken, 13...Bb4
D49.9=Semi-Slaviskt: Meran, Gamla Huvudvarianten, 11.Nxb5 axb5
D49.10=Semi-Slaviskt: Meran, Gamla Huvudvarianten, Botvinnikvarianten
D50.1=Avb�jd damgambit: 4.Bg5
D50.2=Avb�jd damgambit: 4.Bg5 c6
D50.3=Avb�jd damgambit: 4.Bg5 dxc4
D50.4=Avb�jd damgambit: 4.Bg5 Bb4
D50.5=Avb�jd damgambit: Holl�ndsk-Peruvian gambit
D50.6=Avb�jd damgambit: Holl�ndsk-Peruvian, 5.e3
D50.7=Avb�jd damgambit: Semi-Tarrasch, Pillsburyvarianten
D50.8=Avb�jd damgambit: Semi-Tarrasch, Gamla Pillsbury-varianten
D50.9=Avb�jd damgambit: Semi-Tarrasch, Pillsbury, 6.Nxd4
D50.10=Avb�jd damgambit: Semi-Tarrasch, Pillsbury, 6.Nxd4 e5
D50.11=Avb�jd damgambit: Semi-Tarrasch, Pillsbury, Krausevarianten
D50.12=Avb�jd damgambit: Holl�ndsk-Peruvian, 5.cxd5
D50.13=Avb�jd damgambit: Holl�ndsk-Peruvian, Canal (Venice)varianten
D50.14=Avb�jd damgambit: Holl�ndsk-Peruvian, Prinsvarianten
D50.15=Avb�jd damgambit: Holl�ndsk-Peruvian, Prins, 6.Qxd4 Be7 7.e4 Nc6
D50.16=Avb�jd damgambit: Holl�ndsk-Peruvian, Prins, 6.Qxd4 Be7 7.e4 Nc6 8.Qd2
D51.1=Avb�jd damgambit: 4.Bg5 Nbd7
D51.2=Avb�jd damgambit: 4.Bg5 Nbd7 5.Nf3
D51.3=Avb�jd damgambit: 4.Bg5 Nbd7 5.Nf3 c6
D51.4=Avb�jd damgambit: Rochlinvarianten
D51.5=Avb�jd damgambit: Alekhine 4.Bg5 Nbd7 5.Nf3 c6 6.e4
D51.6=Avb�jd damgambit: 4.Bg5 Nbd7 5.e3
D51.7=Avb�jd damgambit: Manhattanvarianten
D51.8=Avb�jd damgambit: 4.Bg5 Nbd7 5.e3 c6
D51.9=Avb�jd damgambit: Capablancas Anti-Cambridge Springs
D51.10=Avb�jd damgambit: 4.Bg5 Nbd7 5.e3 c6 6.cxd5 cxd5
D51.11=Avb�jd damgambit: 4.Bg5 Nbd7 5.e3 c6 6.Qc2
D52.1=Avb�jd damgambit: 4.Bg5 Nbd7 5.e3 c6 6.Nf3
D52.2=Avb�jd damgambit: Cambridge Springs f�rsvar
D52.3=Avb�jd damgambit: Cambridge Springs, Capablancavarianten
D52.4=Avb�jd damgambit: Cambridge Springs, 7.cxd5
D52.5=Avb�jd damgambit: Cambridge Springs, Jugoslaviska varianten
D52.6=Avb�jd damgambit: Cambridge Springs, Jugoslavisk, 8.Qd2
D52.7=Avb�jd damgambit: Cambridge Springs, 7.Nd2
D52.8=Avb�jd damgambit: Cambridge Springs, Rubinsteinvarianten
D52.9=Avb�jd damgambit: Cambridge Springs, Bogoljubowvarianten
D52.10=Avb�jd damgambit: Cambridge Springs, Bogoljubow, 8.Qc2
D52.11=Avb�jd damgambit: Cambridge Springs, 8.Qc2 dxc4
D52.12=Avb�jd damgambit: Cambridge Springs, 8.Qc2 O-O
D52.13=Avb�jd damgambit: Cambridge Springs, Argentinska varianten
D52.14=Avb�jd damgambit: Cambridge Springs, 8.Qc2 O-O 9.Be2
D52.15=Avb�jd damgambit: Cambridge Springs, 8.Qc2 O-O 9.Be2 e5
D53.1=Avb�jd damgambit: 4.Bg5 Be7
D53.2=Avb�jd damgambit: 4.Bg5 Be7 5.cxd5 Nxd5
D53.3=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3
D53.4=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6
D53.5=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bxf6
D53.6=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bxf6 Bxf6
D53.7=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bxf6 Bxf6 7.e3
D53.8=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bh4
D53.9=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bh4 O-O
D53.10=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bh4 O-O 7.Qc2
D53.11=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 h6 6.Bh4 O-O 7.Rc1
D53.12=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 O-O
D53.13=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 O-O 6.Qc2
D53.14=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 O-O 6.Qc2 Nbd7
D53.15=Avb�jd damgambit: 4.Bg5 Be7 5.Nf3 O-O 6.Qc2 c5
D53.16=Avb�jd damgambit: 4.Bg5 Be7 5.e3
D53.17=Avb�jd damgambit: Tidig Lasker variant
D53.18=Avb�jd damgambit: 4.Bg5 Be7 5.e3 Nbd7
D53.19=Avb�jd damgambit: 4.Bg5 Be7 5.e3 Nbd7 6.Nf3
D53.20=Avb�jd damgambit: 4.Bg5 Be7 5.e3 h6
D53.21=Avb�jd damgambit: 4.Bg5 Be7 5.e3 O-O
D53.22=Avb�jd damgambit: 4.Bg5 Be7 5.e3 O-O 6.Qc2
D53.23=Avb�jd damgambit: 4.Bg5 Be7 5.e3 O-O 6.Qc2 c5
D54.1=Avb�jd damgambit: Anti-Neo-Orthodoxvarianten
D54.2=Avb�jd damgambit: Anti-Neo-Orthodoxvarianten
D54.3=Avb�jd damgambit: Anti-Neo-Orthodox, 7.Bh4 b6
D54.4=Avb�jd damgambit: Anti-Neo-Orthodox, 8.cxd5 Nxd5 9.Nxd5
D54.5=Avb�jd damgambit: Anti-Neo-Orthodox, Huvudvarianten
D54.6=Avb�jd damgambit: Anti-Neo-Orthodox, Huvudvarianten, 11.Be2
D55.1=Avb�jd damgambit: 6.Nf3
D55.2=Avb�jd damgambit: Lasker utan ...h6
D55.3=Avb�jd damgambit: 6.Nf3 b6
D55.4=Avb�jd damgambit: 6.Nf3 b6 7.Be2
D55.5=Avb�jd damgambit: 6.Nf3 b6 7.cxd5 exd5
D55.6=Avb�jd damgambit: 6.Nf3 b6 7.cxd5 Nxd5
D55.7=Avb�jd damgambit: Neo-Orthodoxvarianten
D55.8=Avb�jd damgambit: Neo-Orthodox, 7.Bxf6
D55.9=Avb�jd damgambit: Neo-Orthodox, 7.Bxf6 Bxf6 8.Qb3
D55.10=Avb�jd damgambit: Neo-Orthodox, Gligoricvarianten
D55.11=Avb�jd damgambit: Neo-Orthodox, Petrosianvarianten
D56.1=Avb�jd damgambit: Neo-Orthodox, 7.Bh4
D56.2=Avb�jd damgambit: Laskers f�rsvar
D56.3=Avb�jd damgambit: Laskers f�rsvar, 9.Nxe4
D56.4=Avb�jd damgambit: Laskers f�rsvar, Teichmannvarianten
D56.5=Avb�jd damgambit: Laskers f�rsvar, Teichmann, 9...c6
D56.6=Avb�jd damgambit: Laskers f�rsvar, Teichmann, 9...Nxc3
D56.7=Avb�jd damgambit: Laskers f�rsvar, 9.Rc1
D56.8=Avb�jd damgambit: Laskers f�rsvar, 9.Rc1 c6
D56.9=Avb�jd damgambit: Laskers f�rsvar, 9.Rc1 c6 10.Bd3
D57.1=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten
D57.2=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten
D57.3=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten
D57.4=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten, 11.Qb3
D57.5=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten, Bernsteinvarianten
D57.6=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten, Bernstein, 12.c4 dxc4 13.Bxc4
D57.7=Avb�jd damgambit: Laskers f�rsvar, Huvudvarianten, 11.Qb3 Rd8
D58.1=Avb�jd damgambit: Tartakowersystemet
D58.2=Avb�jd damgambit: Tartakower, 8.Qb3
D58.3=Avb�jd damgambit: Tartakower, 8.Qc2
D58.4=Avb�jd damgambit: Tartakower, 8.Bxf6
D58.5=Avb�jd damgambit: Tartakower, 8.Bd3
D58.6=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7
D58.7=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O
D58.8=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7
D58.9=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Bg3
D58.10=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Rc1
D58.11=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Rc1 c5
D58.12=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Qe2
D58.13=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Qe2 c5
D58.14=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Qe2 c5 11.Bg3
D58.15=Avb�jd damgambit: Tartakower, 8.Bd3 Bb7 9.O-O Nbd7 10.Qe2 c5 11.Rfd1
D58.16=Avb�jd damgambit: Tartakower, 8.Be2
D58.17=Avb�jd damgambit: Tartakower, 8.Be2 Bb7
D58.18=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5
D58.19=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5
D58.20=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5 11.O-O
D58.21=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5 11.b4
D58.22=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5 11.b4 c5
D58.23=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5 11.b4 c6
D58.24=Avb�jd damgambit: Tartakower, 8.Be2 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5 11.b4 c6 12.O-O
D58.25=Avb�jd damgambit: Tartakower, 8.Rc1
D58.26=Avb�jd damgambit: Tartakower, 8.Rc1 Bb7
D58.27=Avb�jd damgambit: Tartakower, 8.Rc1 Bb7 9.cxd5
D58.28=Avb�jd damgambit: Tartakower, 8.Rc1 Bb7 9.cxd5 exd5
D58.29=Avb�jd damgambit: Tartakower, 8.Rc1 Bb7 9.Bxf6
D58.30=Avb�jd damgambit: Tartakower, 8.Rc1 Bb7 9.Bxf6 Bxf6 10.cxd5 exd5
D58.31=Avb�jd damgambit: Tartakower, 8.cxd5
D58.32=Avb�jd damgambit: Tartakower, 8.cxd5 exd5
D58.33=Avb�jd damgambit: Tartakower, 8.cxd5 exd5 9.Bd3
D59.1=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5
D59.2=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Nxd5
D59.3=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7
D59.4=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7
D59.5=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1
D59.6=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1 Bb7
D59.7=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1 Bb7 11.Nxd5
D59.8=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1 Bb7 11.Nxd5 Bxd5
D59.9=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1 Bb7 11.Bd3
D59.10=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Rc1 Bb7 11.Be2
D59.11=Avb�jd damgambit: Tartakower, 8.cxd5 Nxd5 9.Bxe7 Qxe7 10.Nxd5
D59.12=Avb�jd damgambit: Tartakower, Huvudvarianten, 11.Rc1
D59.13=Avb�jd damgambit: Tartakower, Huvudvarianten, 11.Rc1
D59.14=Avb�jd damgambit: Tartakower, Huvudvarianten, 11.Rc1 Be6
D59.15=Avb�jd damgambit: Tartakower, Huvudvarianten, 12.Bd3
D59.16=Avb�jd damgambit: Tartakower, Huvudvarianten, 12.Qa4
D59.17=Avb�jd damgambit: Tartakower, Huvudvarianten, 12.Qa4 c5
D60.1=Avb�jd damgambit: Orthodoxt f�rsvar
D60.2=Avb�jd damgambit: Orthodox, 7.cxd5 Nxd5
D60.3=Avb�jd damgambit: Orthodox, Rauzervarianten
D60.4=Avb�jd damgambit: Orthodox, Rauzervarianten
D60.5=Avb�jd damgambit: Orthodox, Botvinnikvarianten
D60.6=Avb�jd damgambit: Orthodox, Botvinnik, 7...b6
D60.7=Avb�jd damgambit: Orthodox, Botvinnik, 7...c6
D60.8=Avb�jd damgambit: Orthodox, Botvinnik, 7...dxc4
D60.9=Avb�jd damgambit: Orthodox, Botvinnik, 7...dxc4 8.Bxc4
D60.10=Avb�jd damgambit: Orthodox, Botvinnik, 8...a6
D60.11=Avb�jd damgambit: Orthodox, Botvinnik, 8...c5
D60.12=Avb�jd damgambit: Orthodox, Botvinnik, 8...c5 9.O-O a6
D61.1=Avb�jd damgambit: Orthodox, Rubinsteinvarianten
D61.2=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 h6
D61.3=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 h6 8.Bh4
D61.4=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 h6 8.Bh4 c5
D61.5=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 a6
D61.6=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c6
D61.7=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c6 8.a3
D61.8=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c6 8.Bd3
D61.9=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c6 8.Bd3 dxc4 9.Bxc4
D61.10=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c6 8.Rd1
D61.11=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5
D61.12=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.Rd1
D61.13=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.O-O-O
D62.1=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5
D62.2=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5 cxd4
D62.3=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5 exd5
D62.4=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5 exd5 9.Bd3
D62.5=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5 Nxd5
D62.6=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5 Nxd5 9.Bxe7 Qxe7
D62.7=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5, Huvudvarianten
D62.8=Avb�jd damgambit: Orthodox, Rubinstein, 7.Qc2 c5 8.cxd5, Huvudvarianten, 11.Bd3
D63.1=Avb�jd damgambit: Orthodox, 7.Rc1
D63.2=Avb�jd damgambit: Orthodox, 7.Rc1 Re8
D63.3=Avb�jd damgambit: Orthodox, 7.Rc1 h6
D63.4=Avb�jd damgambit: Orthodox, 7.Rc1 h6 8.Bh4
D63.5=Avb�jd damgambit: Orthodox, 7.Rc1 dxc4
D63.6=Avb�jd damgambit: Orthodox, 7.Rc1 dxc4 8.Bxc4 a6
D63.7=Avb�jd damgambit: Orthodox, 7.Rc1 b6
D63.8=Avb�jd damgambit: Orthodox, 7.Rc1 b6
D63.9=Avb�jd damgambit: Orthodox, 7.Rc1 b6, Durasvarianten
D63.10=Avb�jd damgambit: Orthodox, 7.Rc1 b6, Pillsburys attack
D63.11=Avb�jd damgambit: Orthodox, 7.Rc1 b6, Capablancavarianten
D63.12=Avb�jd damgambit: Orthodox, Schweiziskvarianten
D63.13=Avb�jd damgambit: Orthodox, Schweizisk, 8.a3
D63.14=Avb�jd damgambit: Orthodox, Schweizisk, 8.c5
D63.15=Avb�jd damgambit: Orthodox, Schweizisk, 8.c5 c6
D63.16=Avb�jd damgambit: Orthodox, Schweizisk, Karlsbadvarianten
D63.17=Avb�jd damgambit: Orthodox, Schweizisk, Karlsbadvarianten
D63.18=Avb�jd damgambit: Orthodox, Schweizisk, Karlsbad, 9.Bd3
D63.19=Avb�jd damgambit: Orthodox, Schweizisk, Karlsbad, 9.Bd3 Re8
D63.20=Avb�jd damgambit: Orthodox, Schweizisk, Karlsbad, 9.Bd3 c6
D63.21=Avb�jd damgambit: Orthodox, 7.Rc1 c6
D63.22=Avb�jd damgambit: Orthodox, 7.Rc1 c6 8.a3
D64.1=Avb�jd damgambit: Orthodox, Rubinsteinattack
D64.2=Avb�jd damgambit: Orthodox, Rubinsteinattack, 8...dxc4
D64.3=Avb�jd damgambit: Orthodox, Rubinsteinattack, Wolfvarianten
D64.4=Avb�jd damgambit: Orthodox, Rubinsteinattack, 8...Re8
D64.5=Avb�jd damgambit: Orthodox, Rubinsteinattack, 8...Re8 9.a3
D64.6=Avb�jd damgambit: Orthodox, Rubinsteinattack, 8...Re8 9.a3 a6
D64.7=Avb�jd damgambit: Orthodox, Rubinsteinattack, 8...h6
D64.8=Avb�jd damgambit: Orthodox, Rubinsteinattack, Carlsbadvarianten
D64.9=Avb�jd damgambit: Orthodox, Rubinsteinattack, Gr�nfeldvarianten
D64.10=Avb�jd damgambit: Orthodox, Rubinsteinattack, Gr�nfeldvarianten, 9...h6
D64.11=Avb�jd damgambit: Orthodox, Rubinsteinattack, Gr�nfeldvarianten, 9...h6 10.Bh4
D65.1=Avb�jd damgambit: Orthodox, Rubinsteinattack, 9.cxd5
D65.2=Avb�jd damgambit: Orthodox, Rubinsteinattack, 9.cxd5 Nxd5
D65.3=Avb�jd damgambit: Orthodox, Rubinsteinattack, 9.cxd5 exd5
D65.4=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 h6
D65.5=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 h6 11.Bh4
D65.6=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 Re8
D65.7=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 Re8 11.O-O Nf8
D65.8=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 Re8 11.O-O Nf8 12.Ne5
D65.9=Avb�jd damgambit: Orthodox, Rubinstein, 9.cxd5 exd5 10.Bd3 Re8 11.O-O Nf8 12.h3
D66.1=Avb�jd damgambit: Orthodox, Huvudvarianten
D66.2=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...a6
D66.3=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...h6
D66.4=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...h6 9.Bh4
D66.5=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...h6 9.Bh4 dxc4
D66.6=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...h6 9.Bh4 dxc4 10.Bxc4
D66.7=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...h6 9.Bh4 dxc4 10.Bxc4 b5
D66.8=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...Re8
D66.9=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...dxc4
D66.10=Avb�jd damgambit: Orthodox, Huvudvarianten, 8...dxc4
D66.11=Avb�jd damgambit: Orthodox, Huvudvarianten, Fianchettovarianten
D66.12=Avb�jd damgambit: Orthodox, Huvudvarianten, Fianchettovarianten
D66.13=Avb�jd damgambit: Orthodox, Huvudvarianten, Fianchetto, 11.O-O
D66.14=Avb�jd damgambit: Orthodox, Huvudvarianten, Fianchetto, 11.e4
D67.1=Avb�jd damgambit: Orthodox, Huvudvarianten, Capablancas befriande man�ver
D67.2=Avb�jd damgambit: Orthodox, Huvudvarianten, Janowskivarianten
D67.3=Avb�jd damgambit: Orthodox, Huvudvarianten, Capablancavarianten
D67.4=Avb�jd damgambit: Orthodox, Huvudvarianten, Alekhinevarianten
D67.5=Avb�jd damgambit: Orthodox, Huvudvarianten, Alekhine, 11...e5 (Lasker)
D67.6=Avb�jd damgambit: Orthodox, Huvudvarianten, Alekhine, 11...N5f6
D67.7=Avb�jd damgambit: Orthodox, Huvudvarianten, Capablanca, 11.O-O
D67.8=Avb�jd damgambit: Orthodox, Huvudvarianten, Capablanca, 11.O-O Nxc3
D68.1=Avb�jd damgambit: Orthodox, Klassiska varianten
D68.2=Avb�jd damgambit: Orthodox, Klassisk, 13.Bb3
D68.3=Avb�jd damgambit: Orthodox, Klassisk, Maroczyvarianten
D68.4=Avb�jd damgambit: Orthodox, Klassisk, Maroczy, 13...exd4
D68.5=Avb�jd damgambit: Orthodox, Klassisk, Vidmarvarianten
D68.6=Avb�jd damgambit: Orthodox, Klassisk, Vidmar, 13...e4
D68.7=Avb�jd damgambit: Orthodox, Klassisk, Vidmar, 13...exd4
D68.8=Avb�jd damgambit: Orthodox, Klassisk, Vidmar, 13...exd4 14.exd4 Nb6
D69.1=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5
D69.2=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5
D69.3=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5: 15.f4
D69.4=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5: 15.f4 Qe4
D69.5=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5: 15.f4 Qf6
D69.6=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5: 15.f4 Qf6 16.f5
D69.7=Avb�jd damgambit: Orthodox, Klassisk, 13.dxe5: 15.f4 Qf6 16.e4
D70.1=Neo-Gr�nfeld: 3.Nf3 d5
D70.2=Neo-Gr�nfeld: Alekhines Anti-Gr�nfeld
D70.3=Neo-Gr�nfeld: Alekhines, 5.e4 Nb6
D70.4=Neo-Gr�nfeld: Alekhines, 7.Be3 O-O
D70.5=Neo-Gr�nfeld: 3.g3 d5
D70.6=Neo-Gr�nfeld: 4.cxd5
D70.7=Neo-Gr�nfeld: 4.Bg2
D70.8=Neo-Gr�nfeld: 4.Bg2 c6
D70.9=Neo-Gr�nfeld: 4.Bg2 Bg7
D71.1=Neo-Gr�nfeld, 5.cxd5 Nxd5
D71.2=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.Nc3
D71.3=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.Nc3 Nxc3
D71.4=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.Nc3 Nxc3 7.bxc3 c5
D71.5=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.Nc3 Nb6
D71.6=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4
D71.7=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6
D71.8=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb4
D71.9=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb4 7.d5
D72.1=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2
D72.2=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2 Nc6
D72.3=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2 e5
D72.4=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2 c5
D72.5=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2 O-O
D72.6=Neo-Gr�nfeld, 5.cxd5 Nxd5 6.e4 Nb6 7.Ne2 O-O 8.O-O
D73.1=Neo-Gr�nfeld, 5.Nf3
D73.2=Neo-Gr�nfeld, 5.Nf3 c6
D73.3=Neo-Gr�nfeld, 5.Nf3 c6 6.cxd5
D73.4=Neo-Gr�nfeld, 5.Nf3 c6 6.cxd5 cxd5
D73.5=Neo-Gr�nfeld, 5.Nf3 c6 6.cxd5 cxd5 7.Nc3
D73.6=Neo-Gr�nfeld, 5.Nf3 c5
D73.7=Neo-Gr�nfeld, 5.Nf3 dxc4
D73.8=Neo-Gr�nfeld, 5.Nf3 dxc4 6.Na3
D73.9=Neo-Gr�nfeld, 5.Nf3 O-O
D73.10=Neo-Gr�nfeld, 6.Qb3
D73.11=Neo-Gr�nfeld, 6.Nc3
D73.12=Neo-Gr�nfeld, 6.cxd5
D73.13=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.e4
D74.1=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O
D74.2=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Na6
D74.3=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nc6
D74.4=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c6
D74.5=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5
D74.6=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.e4
D74.7=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.e4 Nf6
D74.8=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.e4 Nf6 9.e5 Nd5
D75.1=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.Nc3
D75.2=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.Nc3 Nxc3
D75.3=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.Nc3 Nxc3 9.bxc3 cxd4
D75.4=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.dxc5
D75.5=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O c5 8.dxc5 Na6
D76.1=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6
D76.2=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3
D76.3=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6
D76.4=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.e3
D76.5=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.e3 e5
D76.6=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.e3 Re8
D76.7=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.d5
D76.8=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.d5 Na5
D76.9=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.d5 Na5 10.e4
D76.10=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.d5 Na5 10.e4 c6
D76.11=Neo-Gr�nfeld, 6.cxd5 Nxd5 7.O-O Nb6 8.Nc3 Nc6 9.d5 Na5 10.e4 c6 11.Bg5
D77.1=Neo-Gr�nfeld, 6.O-O
D77.2=Neo-Gr�nfeld, 6.O-O e6
D77.3=Neo-Gr�nfeld, 6.O-O c5
D77.4=Neo-Gr�nfeld, 6.O-O c5 7.dxc5 dxc4
D77.5=Neo-Gr�nfeld, 6.O-O dxc4
D77.6=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3
D77.7=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Na6
D77.8=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 c3
D77.9=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 c3 8.bxc3 c5
D77.10=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 c3 8.bxc3 c5 9.e3
D77.11=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Nc6
D77.12=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Nc6 8.Nxc4
D77.13=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Nc6 8.Nxc4 Be6
D77.14=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Nc6 8.Nxc4 Be6 9.b3
D77.15=Neo-Gr�nfeld, 6.O-O dxc4 7.Na3 Nc6 8.Nxc4 Be6 9.b3 Bd5
D78.1=Neo-Gr�nfeld, 6.O-O c6
D78.2=Neo-Gr�nfeld, 6.O-O c6 7.Na3
D78.8=Neo-Gr�nfeld, 6.O-O c6 7.Ne5
D78.3=Neo-Gr�nfeld, 6.O-O c6 7.Qa4
D78.9=Neo-Gr�nfeld, 6.O-O c6 7.Nc3
D78.10=Neo-Gr�nfeld, 6.O-O c6 7.Nc3 dxc4
D78.4=Neo-Gr�nfeld, 6.O-O c6 7.Qb3
D78.5=Neo-Gr�nfeld, 6.O-O c6 7.Qb3 Qb6
D78.6=Neo-Gr�nfeld, 6.O-O c6 7.Qb3 dxc4
D78.7=Neo-Gr�nfeld, 6.O-O c6 7.Qb3 dxc4
D78.11=Neo-Gr�nfeld, 6.O-O c6 7.Nbd2
D78.12=Neo-Gr�nfeld, 6.O-O c6 7.Nbd2 Nbd7
D78.13=Neo-Gr�nfeld, 6.O-O c6 7.Nbd2 Ne4
D78.14=Neo-Gr�nfeld, 6.O-O c6 7.Nbd2 Bf5
D78.15=Neo-Gr�nfeld, 6.O-O c6 7.b3
D78.16=Neo-Gr�nfeld, 6.O-O c6 7.b3 Bf5
D78.17=Neo-Gr�nfeld, 6.O-O c6 7.b3 Ne4
D79.1=Neo-Gr�nfeld, 6.O-O c6 7.cxd5
D79.2=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5
D79.3=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3
D79.4=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 e6
D79.5=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Ne4
D79.6=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Ne4 9.Ne5
D79.7=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Ne4 9.Nxe4
D79.8=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Nc6
D79.9=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Nc6 9.Ne5
D79.10=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Nc3 Nc6 9.Ne5 e6
D79.11=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Ne5
D79.12=Neo-Gr�nfeld, 6.O-O c6 7.cxd5 cxd5 8.Ne5 e6
D79.13=Neo-Gr�nfeld, Huvudvarianten
D79.14=Neo-Gr�nfeld, Huvudvarianten, 10.f4
D79.15=Neo-Gr�nfeld, Huvudvarianten, 10.f4 Nc6
D79.16=Neo-Gr�nfeld, Huvudvarianten, 10.f4 Nc6 11.Be3
D79.17=Neo-Gr�nfeld, Huvudvarianten, 10.f4 Nc6 11.Be3 f6
D79.18=Neo-Gr�nfeld, Huvudvarianten, 10.f4 Nc6 11.Be3 Nb6
D79.19=Neo-Gr�nfeld, Huvudvarianten, 10.f4 Nc6 11.Be3 Nb6 12.Bf2
D80.1=Gr�nfelds f�rsvar
D80.2=Gr�nfeld: Tagg/Gibbon gambit
D80.3=Gr�nfeld: 4.h4
D80.4=Gr�nfeld: 4.g3
D80.5=Gr�nfeld: 4.f3
D80.6=Gr�nfeld: 4.e3
D80.7=Gr�nfeld: 4.e3 Bg7
D80.8=Gr�nfeld: 4.e3 Bg7 5.Qb3
D80.9=Gr�nfeld: Stockholmvarianten
D80.10=Gr�nfeld: Stockholm, 4...Ne4
D80.11=Gr�nfeld: Stockholm, 4...Ne4 5.Nxe4
D80.12=Gr�nfeld: Stockholm, Lundinvarianten
D80.13=Gr�nfeld: Stockholm, 4...Ne4 5.Bf4
D80.14=Gr�nfeld: Stockholm, Taimanovvarianten
D80.15=Gr�nfeld: Stockholm, Taimanov, 5...Nxc3
D80.16=Gr�nfeld: Stockholm, Taimanov, 5...Nxc3 6.bxc3 Bg7
D81.1=Gr�nfeld: Tidiga ryska varianten
D81.2=Gr�nfeld: Tidiga ryska varianten
D81.3=Gr�nfeld: Tidig rysk, 5...Be6
D81.4=Gr�nfeld: Tidig rysk, 5...Be6 6.Qb5+
D81.5=Gr�nfeld: Tidig rysk, Adorjan gambit
D81.6=Gr�nfeld: Tidig rysk, 5...Bg7
D81.7=Gr�nfeld: Tidig rysk, 5...Bg7 6.e4
D81.8=Gr�nfeld: Tidig rysk, 5...Bg7 6.e4 O-O
D82.1=Gr�nfeld: 4.Bf4
D82.2=Gr�nfeld: 4.Bf4 Bg7
D82.3=Gr�nfeld: 4.Bf4 Bg7 5.e3
D82.4=Gr�nfeld: 4.Bf4 Bg7 5.e3 c5
D82.5=Gr�nfeld: 4.Bf4 Bg7 5.e3 c5 6.dxc5 Qa5
D82.6=Gr�nfeld: 4.Bf4 Bg7 5.e3 c5 6.dxc5 Qa5 7.Qa4+
D82.7=Gr�nfeld: 4.Bf4 Bg7 5.e3 c5 6.dxc5 Qa5 7.Rc1
D83.1=Gr�nfeld: Gr�nfeld gambit
D83.2=Gr�nfeld: Gr�nfeld gambit, 6.Qb3
D83.3=Gr�nfeld: Gr�nfeld gambit, Capablancavarianten
D83.4=Gr�nfeld: Gr�nfeld gambit, Capablancavarianten
D83.5=Gr�nfeld: Gr�nfeld gambit, Botvinnikvarianten
D84.1=Gr�nfeld: Antagen Gr�nfeldgambit
D84.2=Gr�nfeld: Antagen Gr�nfeldgambit
D84.3=Gr�nfeld: Antagen Gr�nfeldgambit, 8...b6
D84.4=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Bf5
D84.5=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Na6
D84.6=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Na6 9.Bxa6 Qxg2
D84.7=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Nc6
D84.8=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Nc6 9.Ne2
D84.9=Gr�nfeld: Antagen Gr�nfeldgambit, 8...Nc6 9.Ne2 Bg4
D85.1=Gr�nfeld: Avbytesvarianten
D85.2=Gr�nfeld: Avbytesvarianten
D85.3=Gr�nfeld: Avbyte, 5.g3
D85.4=Gr�nfeld: Avbyte, 5.Na4
D85.5=Gr�nfeld: Avbyte, 5.Bd2
D85.6=Gr�nfeld: Avbyte, 5.Bd2 Bg7 6.e4 Nb6
D85.7=Gr�nfeld: Avbyte, 5.Bd2 Bg7 6.e4 Nb6 7.Be3
D85.8=Gr�nfeld: Avbyte, 5.e4
D85.9=Gr�nfeld: Avbyte, 5.e4 Nb6
D85.10=Gr�nfeld: Avbyte, 5.e4 Nxc3
D85.11=Gr�nfeld: Avbyte, 5.e4 Nxc3 6.bxc3 c5
D85.12=Gr�nfeld: Avbyte, 5.e4 Nxc3 6.bxc3 Bg7
D85.13=Gr�nfeld: Avbyte, 7.Ba3
D85.14=Gr�nfeld: Avbyte, 7.Bb5+
D85.15=Gr�nfeld: Avbyte, 7.Bb5+ c6
D85.16=Gr�nfeld: Avbyte, 7.Bb5+ c6 8.Ba4
D85.17=Gr�nfeld: Avbyte, 7.Bb5+ c6 8.Ba4 O-O
D85.18=Gr�nfeld: Avbyte, 7.Be3
D85.19=Gr�nfeld: Avbyte, 7.Be3 c5
D85.20=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2
D85.21=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 O-O
D85.22=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 O-O 9.Rc1
D85.23=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 Qa5
D85.24=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 Qa5 9.Rc1
D85.25=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 Qa5 9.Rb1
D85.26=Gr�nfeld: Avbyte, 7.Be3 c5 8.Qd2 Qa5 9.Rb1 b6
D85.27=Gr�nfeld: Modernt avbyte
D85.28=Gr�nfeld: Modernt avbyte, 7...O-O
D85.29=Gr�nfeld: Modernt avbyte, 7...c5
D85.30=Gr�nfeld: Modernt avbyte, 8.Bb5+
D85.31=Gr�nfeld: Modernt avbyte, 8.Be2
D85.32=Gr�nfeld: Modernt avbyte, 8.Be2 O-O
D85.33=Gr�nfeld: Modernt avbyte, 8.Be2 O-O 9.O-O
D85.34=Gr�nfeld: Modernt avbyte, 8.Be2 O-O 9.O-O b6
D85.35=Gr�nfeld: Modernt avbyte, 8.Be2 O-O 9.O-O Nc6
D85.36=Gr�nfeld: Modernt avbyte, 8.Rb1
D85.37=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O
D85.38=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2
D85.39=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 Qa5
D85.40=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 b6
D85.41=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 Nc6
D85.42=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 Nc6, Huvudvarianten
D85.43=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 Nc6, Huvudvarianten, 12...e6
D85.44=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 cd
D85.45=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 cd 10.cd
D85.46=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 cd 10.cd Qa5+
D85.47=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 cd 10.cd Qa5+ 11.Qd2
D85.48=Gr�nfeld: Modernt avbyte, 8.Rb1 O-O 9.Be2 cd 10.cd Qa5+ 11.Bd2
D85.49=Gr�nfeld: Modernt avbyte, 8.Rb1, 10...Qa5+ 11.Bd2 Qxa2 12.O-O Bg4
D85.50=Gr�nfeld: Modernt avbyte, 8.Rb1, 10...Qa5+ 11.Bd2 Qxa2 12.O-O Bg4 13.Bg5
D85.51=Gr�nfeld: Modernt avbyte, 8.Be3
D85.52=Gr�nfeld: Modernt avbyte, 8.Be3 Bg4
D85.53=Gr�nfeld: Modernt avbyte, 8.Be3 Nc6
D85.54=Gr�nfeld: Modernt avbyte, 8.Be3 Qa5
D85.55=Gr�nfeld: Modernt avbyte, 8.Be3 Qa5 9.Qd2
D85.56=Gr�nfeld: Modernt avbyte, 8.Be3 Qa5 9.Qd2 Nc6 10.Rc1
D85.57=Gr�nfeld: Modernt avbyte, 8.Be3 O-O
D85.58=Gr�nfeld: Modernt avbyte, 8.Be3 O-O 9.Rc1 Qa5
D85.59=Gr�nfeld: Modernt avbyte, 8.Be3 O-O 9.Rc1 Qa5 10.Qd2
D85.60=Gr�nfeld: Modernt avbyte, 8.Be3 O-O 9.Rc1 Qa5 Dambyte, 12.Kxd2
D85.61=Gr�nfeld: Modernt avbyte, 8.Be3 O-O 9.Rc1 Qa5 Dambyte, 12.Nxd2
D86.1=Gr�nfeld: Klassiskt avbyte
D86.2=Gr�nfeld: Klassiskt avbyte, 7...b6
D86.3=Gr�nfeld: Klassiskt avbyte, 7...c5
D86.4=Gr�nfeld: Klassiskt avbyte, 7...O-O
D86.5=Gr�nfeld: Klassiskt avbyte, 8.Ne2
D86.6=Gr�nfeld: Klassiskt avbyte, Larsenvarianten
D86.7=Gr�nfeld: Klassiskt avbyte, Simagin
D86.8=Gr�nfeld: Klassiskt avbyte, Simagin, 9.h4
D86.9=Gr�nfeld: Klassiskt avbyte, Simagin, 9.O-O
D86.10=Gr�nfeld: Klassiskt avbyte, Simagin F�rb�ttrad
D86.11=Gr�nfeld: Klassiskt avbyte, Simagin F�rb�ttrad, 9.Be3
D86.12=Gr�nfeld: Klassiskt avbyte, Simagin F�rb�ttrad, 9.O-O
D86.13=Gr�nfeld: Klassiskt avbyte, Simagin F�rb�ttrad, 9.O-O e5
D86.14=Gr�nfeld: Klassiskt avbyte, Simagin F�rb�ttrad, 9.O-O b6
D87.1=Gr�nfeld: Klassiskt avbyte, 8...c5
D87.2=Gr�nfeld: Klassiskt avbyte, 8...c5 9.Be3
D87.3=Gr�nfeld: Klassiskt avbyte, 8...c5 9.Be3 Qa5
D87.4=Gr�nfeld: Klassiskt avbyte, 8...c5 9.Be3 Qa5
D87.5=Gr�nfeld: Klassiskt avbyte, 8...c5 9.Be3 Nc6
D87.6=Gr�nfeld: Klassiskt avbyte, 9.O-O
D87.7=Gr�nfeld: Klassiskt avbyte, 9.O-O Nc6
D87.8=Gr�nfeld: Klassiskt avbyte, 9.O-O Nc6 10.Be3
D87.9=Gr�nfeld: Klassiskt avbyte, 10.Be3 Qa5
D87.10=Gr�nfeld: Klassiskt avbyte, 10.Be3 Na5
D87.11=Gr�nfeld: Klassiskt avbyte, 10.Be3 Qc7
D87.12=Gr�nfeld: Klassiskt avbyte, 10.Be3 Qc7 11.Rc1 Rd8
D87.13=Gr�nfeld: Klassiskt avbyte, 10.Be3 Qc7 11.Rc1 Rd8 12.Qd2
D87.14=Gr�nfeld: Klassiskt avbyte, 10.Be3 Qc7 11.Rc1 Rd8 12.Bf4
D87.15=Gr�nfeld: Klassiskt avbyte, 10.Be3 Bg4
D87.16=Gr�nfeld: Klassiskt avbyte, 10.Be3 Bg4 11.f3 Na5 12.Bd5
D87.17=Gr�nfeld: Klassiskt avbyte, Sevillevarianten
D88.1=Gr�nfeld: Klassiskt avbyte, Huvudvarianten
D88.2=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4
D88.3=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Na5
D88.4=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Na5 12.Bd3
D88.5=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Bg4
D88.6=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Bg4 12.f3
D88.7=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Bg4 12.f3 Na5
D88.8=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, Neo-Seville
D88.9=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 11.cxd4 Bg4 12.f3 Na5 13.Bd5
D89.1=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 13.Bd3
D89.2=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 13.Bd3 Be6
D89.3=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, 13.Bd3 Be6 14.Rc1
D89.4=Gr�nfeld: Klassiskt avbyte, 14.Rc1 Bxa2 15.Qa4 Be6 16.d5 Be7 17.Qb4
D89.5=Gr�nfeld: Klassiskt avbyte, 14.Rc1 Bxa2 15.Qa4 med 17.Qb4 b6
D89.6=Gr�nfeld: Klassiskt avbyte, 14.Rc1 Bxa2 15.Qa4 med 17.Qb4 e6
D89.7=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, Sokolskyvarianten
D89.8=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, Sokolsky, 16.Rb1
D89.9=Gr�nfeld: Klassiskt avbyte, Huvudvarianten, Sokolsky, 16.Bh6
D90.1=Gr�nfeld: Trespringarvarianten
D90.2=Gr�nfeld: Schlechtervarianten
D90.3=Gr�nfeld: Schlechter, 5.Qb3
D90.4=Gr�nfeld: Schlechter, Avbyte
D90.5=Gr�nfeld: Schlechter, Avbyte
D90.6=Gr�nfeld: Trespringarvarianten
D90.7=Gr�nfeld: Trespringar, 5.g3
D90.8=Gr�nfeld: Flohrvarianten
D90.9=Gr�nfeld: Trespringaravbyte
D90.10=Gr�nfeld: Trespringaravbyte
D90.11=Gr�nfeld: Trespringaravbyte, Romanishinvarianten
D90.12=Gr�nfeld: Trespringaravbyte, 6.Bd2
D90.13=Gr�nfeld: Trespringaravbyte, 6.Bd2 O-O
D90.14=Gr�nfeld: Trespringaravbyte, 6.Bd2 O-O 7.Rc1
D91.1=Gr�nfeld: 5.Bg5
D91.2=Gr�nfeld: 5.Bg5 c6
D91.3=Gr�nfeld: 5.Bg5 dxc4
D91.4=Gr�nfeld: 5.Bg5 dxc4 6.e4
D91.5=Gr�nfeld: 5.Bg5 Ne4
D91.6=Gr�nfeld: 5.Bg5 Ne4 6.Bf4
D91.7=Gr�nfeld: 5.Bg5 Ne4 6.Bh4
D91.8=Gr�nfeld: 5.Bg5 Ne4 6.Bh4 Nxc3
D91.9=Gr�nfeld: 5.Bg5 Ne4 6.Bh4 Nxc3 7.bxc3 dxc4
D91.10=Gr�nfeld: 5.Bg5 Ne4 6.cxd5
D91.11=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5
D91.12=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 c6
D91.13=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6
D91.14=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Qd2
D91.15=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Qd2 exd5
D91.16=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Qd2 exd5: 11.h4 h6
D91.17=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3
D91.18=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3
D91.19=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O
D91.20=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.Bd3
D91.21=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.Bd3
D91.22=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.Be2
D91.23=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.Be2
D91.24=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.b4
D91.25=Gr�nfeld: 5.Bg5 Ne4 6.cxd5 Nxg5 7.Nxg5 e6 8.Nf3 exd5 9.e3 O-O 10.b4 c6
D92.1=Gr�nfeld: 5.Bf4
D92.2=Gr�nfeld: 5.Bf4 c6
D92.3=Gr�nfeld: 5.Bf4 O-O
D92.4=Gr�nfeld: 5.Bf4 O-O 6.Rc1
D92.5=Gr�nfeld: 5.Bf4 O-O 6.Rc1 dxc4
D92.6=Gr�nfeld: 5.Bf4 O-O 6.Rc1 c5
D93.1=Gr�nfeld: 5.Bf4 O-O 6.e3
D93.2=Gr�nfeld: 5.Bf4 O-O 6.e3 c5
D93.3=Gr�nfeld: 5.Bf4 O-O 6.e3 c5 7.dxc5
D93.4=Gr�nfeld: 5.Bf4 O-O 6.e3 c5 7.dxc5 Qa5
D93.5=Gr�nfeld: 5.Bf4 O-O 6.e3 c5 7.dxc5 Qa5 8.Rc1
D93.6=Gr�nfeld: 5.Bf4 O-O 6.e3 c5 7.dxc5 Qa5 8.Rc1 dxc4 9.Bxc4
D93.7=Gr�nfeld: 5.Bf4 O-O 6.e3 c6
D93.8=Gr�nfeld: 5.Bf4 O-O 6.e3 c6 7.Qb3
D93.9=Gr�nfeld: 5.Bf4 O-O 6.e3 c6 7.Rc1
D94.1=Gr�nfeld: 5.e3
D94.2=Gr�nfeld: Slaviskt/Schlecter
D94.3=Gr�nfeld: Slaviskt/Schlecter, 6.Bd3
D94.4=Gr�nfeld: Slaviskt/Schlecter, 6.Be2
D94.5=Gr�nfeld: Slaviskt/Schlecter, 6.Be2 O-O
D94.6=Gr�nfeld: Slaviskt/Schlecter, 6.Be2 O-O 7.O-O
D94.7=Gr�nfeld: 5.e3 O-O
D94.8=Gr�nfeld: Makogonovvarianten
D94.9=Gr�nfeld: Opovcenskyvarianten
D94.10=Gr�nfeld: 5.e3 O-O 6.Be2
D94.11=Gr�nfeld: 5.e3 O-O 6.Be2 c5
D94.12=Gr�nfeld: 5.e3 O-O 6.Bd3
D94.13=Gr�nfeld: 5.e3 O-O 6.Bd3 c6
D94.14=Gr�nfeld: Smyslovs f�rsvar
D94.15=Gr�nfeld: Flohrs f�rsvar
D94.16=Gr�nfeld: 5.e3 O-O 6.cxd5
D94.17=Gr�nfeld: 5.e3 O-O 6.cxd5
D94.18=Gr�nfeld: 5.e3 O-O 6.cxd5 Nxd5 7.Bc4
D95.1=Gr�nfeld: 5.e3 O-O 6.Qb3
D95.2=Gr�nfeld: 5.e3 O-O 6.Qb3 b6
D95.3=Gr�nfeld: 5.e3 O-O 6.Qb3 c6
D95.4=Gr�nfeld: 5.e3 O-O 6.Qb3 c6 7.Bd2 e6
D95.5=Gr�nfeld: 5.e3 O-O 6.Qb3 c6 7.Bd2 e6 8.Bd3
D95.6=Gr�nfeld: Botvinnikvarianten
D95.7=Gr�nfeld: Botvinnik, 7.Bd2
D95.8=Gr�nfeld: 5.e3 O-O 6.Qb3 dxc4
D95.9=Gr�nfeld: 5.e3 O-O 6.Qb3 dxc4 7.Bxc4
D95.10=Gr�nfeld: Pachmanvarianten
D96.1=Gr�nfeld: Ryskta varianten
D96.2=Gr�nfeld: Ryskt, 5...c6
D96.3=Gr�nfeld: Ryskt, 5...c6 6.Bf4
D96.4=Gr�nfeld: Ryskt, 5...c6 6.cxd5 cxd5
D96.5=Gr�nfeld: Ryskt, 5...c6 6.cxd5 Nxd5
D96.6=Gr�nfeld: Ryskt, 5...dxc4
D96.7=Gr�nfeld: Ryskt, 5...dxc4
D96.8=Gr�nfeld: Ryskt, 6...O-O
D96.9=Gr�nfeld: Ryskt, 6...a6
D96.10=Gr�nfeld: Ryskt, 7.Bf4
D96.11=Gr�nfeld: Ryskt, 7.Bf4 c6
D97.1=Gr�nfeld: Ryskt, 7.e4
D97.2=Gr�nfeld: Ryskt, 7.e4 Nfd7
D97.3=Gr�nfeld: Ryskt, Levenfishvarianten
D97.4=Gr�nfeld: Ryskt, Szabovarianten
D97.5=Gr�nfeld: Ryskt, Szabo, 8.Be2
D97.6=Gr�nfeld: Ryskt, Alekhine (Ungersk) variant
D97.7=Gr�nfeld: Ryskt, Alekhine, 8.Be2
D97.8=Gr�nfeld: Ryskt, Alekhine, 8.Be2 b5 9.Qb3
D97.9=Gr�nfeld: Ryskt, Alekhine, 8.Qb3
D97.10=Gr�nfeld: Ryskt, Alekhine, 8.e5
D97.11=Gr�nfeld: Ryskt, Alekhine, 8.e5 b5 9.Qb3
D97.12=Gr�nfeld: Ryskt, Alekhine, 8.e5 b5 9.Qb3 Nfd7
D97.13=Gr�nfeld: Ryskt, Alekhine, 8.e5 b5 9.Qb3 Nfd7 10.Be3
D97.14=Gr�nfeld: Ryskt, Simaginvarianten
D97.15=Gr�nfeld: Ryskt, Simagin, 8.Be2
D97.16=Gr�nfeld: Ryskt, Prinsvarianten
D97.17=Gr�nfeld: Ryskt, Prins, 8.Bf4
D97.18=Gr�nfeld: Ryskt, Prins, 8.Be2
D97.19=Gr�nfeld: Ryskt, Prins, 8.Be2, Huvudvarianten
D98.1=Gr�nfeld: Ryskt, Smyslovvarianten
D98.2=Gr�nfeld: Ryskt, Smyslov, 8.Be2
D98.3=Gr�nfeld: Ryskt, Smyslov, 8.Be2 Nc6
D98.4=Gr�nfeld: Ryskt, Smyslov, 8.Be2 Nc6 9.d5
D98.5=Gr�nfeld: Ryskt, Smyslov, 8.Be3
D98.6=Gr�nfeld: Ryskt, Smyslov, 8.Be3 Nfd7
D98.7=Gr�nfeld: Ryskt, Smyslov, 8.Be3 Nfd7 9.Be2
D98.8=Gr�nfeld: Ryskt, Smyslov, Keresvarianten
D98.9=Gr�nfeld: Ryskt, Smyslov, 8.Be3 Nfd7 9.O-O-O
D98.10=Gr�nfeld: Ryskt, Smyslov, 8.Be3 Nfd7 9.Rd1
D98.11=Gr�nfeld: Ryskt, Smyslov, 8.Be3 Nfd7 9.Rd1 Nc6
D99.1=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten
D99.2=Gr�nfeld: Ryskt, Smyslov, Jugoslavisk
D99.3=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten, 9...Nb6
D99.4=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten, 9...Nb6 10.Rd1
D99.5=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten, 9...Nb6 10.Rd1 e6
D99.6=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten, 9...Nb6 10.Rd1 Nc6
D99.7=Gr�nfeld: Ryskt, Smyslov, Huvudvarianten, 9...Nb6 10.Rd1 Nc6 11.d5 Ne5
E00.1=Dambonde: Neoindiskt
E00.2=Dambonde: Neoindiskt, Devins gambit
E00.3=Dambonde: Anti-Nimzo-Indiskt
E00.4=Dambonde: Anti-Nimzo-Indiskt, 3...d5
E00.5=Neoindisk (Seirawan) attack
E00.6=Dambonde: Neoindiskt
E00.7=Dambonde: Neoindiskt, 3...b6
E00.8=Dambonde: Neoindiskt, 3...b6
E00.9=Dambonde: Neoindiskt, 3...c5
E00.10=Katalansk
E00.11=Katalanskt: Ungersk gambit
E00.12=Katalanskt: 3...c6
E00.13=Katalanskt: 3...c5
E00.14=Katalanskt: 3...c5 4.Nf3
E00.15=Katalanskt: 3...Bb4+
E00.16=Katalanskt: 3...Bb4+ 4.Nd2
E00.17=Katalanskt: 3...Bb4+ 4.Bd2
E00.18=Katalanskt: 3...Bb4+ 4.Bd2 Bxd2+
E00.19=Katalanskt: 3...Bb4+ 4.Bd2 Be7
E00.20=Katalanskt: 3...Bb4+ 4.Bd2 Qe7
E00.21=Katalanskt: 3...Bb4+ 4.Bd2 Qe7
E00.22=Katalanskt: 3...d5
E00.23=Katalanskt: 4.Nf3
E00.24=Katalanskt: 4.Nf3 c6
E00.25=Katalanskt: 4.Nf3 c5
E00.26=Katalanskt: 4.Nf3 Bb4+
E00.27=Katalanskt: 4.Nf3 Bb4+ 5.Bd2
E00.28=Katalanskt: 4.Nf3 Be7
E00.29=Katalanskt: 4.Nf3 dxc4
E00.30=Katalanskt: 4.Nf3 dxc4 5.Qa4+
E00.31=Katalanskt: 4.Nf3 dxc4 5.Qa4+ Nbd7
E01.1=Katalanskt: 4.Bg2
E01.2=Katalanskt: 4...Bb4+
E01.3=Katalanskt: 4...Bb4+ 5.Bd2
E01.4=Katalanskt: 4...Bb4+ 5.Nd2
E01.5=Katalanskt: 4...Bb4+ 5.Nd2 O-O
E01.6=Katalanskt: 4...c6
E01.7=Katalanskt: 4...c6 5.Qc2
E01.8=Katalanskt: 4...c6 5.Nf3
E01.9=Katalanskt: 4...c6 5.Nf3 Nbd7
E01.10=Katalanskt: 4...c5
E01.11=Katalanskt: 4...c5 5.Nf3
E01.12=Katalanskt: �ppet
E02.1=Katalanskt: �ppet, 5.Qa4+
E02.2=Katalanskt: �ppet, 5.Qa4+ Bd7
E02.3=Katalanskt: �ppet, 5.Qa4+ Bd7 6.Qxc4
E02.4=Katalanskt: �ppet, 5.Qa4+ Nbd7
E02.5=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Nf3
E02.6=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Nf3 a6
E02.7=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Nf3 a6 7.Nc3
E03.1=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4
E03.2=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 a6
E03.3=Katalanskt: �ppet, Alekhinevarianten
E03.4=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 a6 7.Nf3
E03.5=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 a6 7.Nf3 b5
E03.6=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 a6 7.Nf3 b5 8.Qc2
E03.7=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 a6 7.Nf3 b5 8.Qc6
E03.8=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5
E03.9=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5 7.Nf3
E03.10=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5 7.Nf3 a6
E03.11=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5 7.Nf3 a6 8.O-O
E03.12=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5 7.Nf3 a6 8.Qc2
E03.13=Katalanskt: �ppet, 5.Qa4+ Nbd7 6.Qxc4 c5 7.Nf3 a6 8.Qc2 b6
E04.1=Katalanskt: �ppet, 5.Nf3
E04.2=Katalanskt: �ppet, 5.Nf3 Bd7
E04.3=Katalanskt: �ppet, 5.Nf3 Bb4+
E04.4=Katalanskt: �ppet, 5.Nf3 Nbd7
E04.5=Katalanskt: �ppet, 5.Nf3 b5
E04.6=Katalanskt: �ppet, 5.Nf3 a6
E04.7=Katalanskt: �ppet, 5.Nf3 a6 6.O-O
E04.8=Katalanskt: �ppet, 5.Nf3 a6 6.O-O b5
E04.9=Katalanskt: �ppet, 5.Nf3 a6 6.O-O b5 7.Ne5
E04.10=Katalanskt: �ppet, 5.Nf3 a6 6.O-O b5 7.Ne5 Nd5 8.a4
E04.11=Katalanskt: �ppet, 5.Nf3 a6 6.O-O Nc6
E04.12=Katalanskt: �ppet, 5.Nf3 a6 6.O-O Nc6 7.e3
E04.13=Katalanskt: �ppet, 5.Nf3 c5
E04.14=Katalanskt: �ppet, 5.Nf3 c5 6.O-O
E04.15=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6
E04.16=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Ne5
E04.17=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Ne5 Bd7 8.Na3
E04.18=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Ne5 Bd7 8.Na3
E04.19=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Qa4
E04.20=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Qa4 cxd4
E04.21=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Qa4 Bd7
E04.22=Katalanskt: �ppet, 5.Nf3 c5 6.O-O Nc6 7.Qa4 Bd7 8.Qxc4
E04.23=Katalanskt: �ppet, 5.Nf3 Nc6
E04.24=Katalanskt: �ppet, 5.Nf3 Nc6 6.O-O
E04.25=Katalanskt: �ppet, 5.Nf3 Nc6 6.O-O Rb8
E04.26=Katalanskt: �ppet, 5.Nf3 Nc6 6.O-O Rb8 7.Nc3
E04.27=Katalanskt: �ppet, 5.Nf3 Nc6 6.Qa4
E04.28=Katalanskt: �ppet, 5.Nf3 Nc6 6.Qa4 Bb4+
E04.29=Katalanskt: �ppet, 5.Nf3 Nc6 6.Qa4 Bb4+ 7.Bd2 Nd5
E05.1=Katalanskt: �ppet, Klassisk
E05.2=Katalanskt: �ppet, Klassisk, 6.Nc3
E05.3=Katalanskt: �ppet, Klassisk, 6.Nc3 O-O
E05.4=Katalanskt: �ppet, Klassisk, 6.Nc3 O-O 7.Ne5
E05.5=Katalanskt: �ppet, Klassisk, 6.O-O
E05.6=Katalanskt: �ppet, Klassisk, 6.O-O O-O
E05.7=Katalanskt: �ppet, Klassisk, 7.Ne5
E05.8=Katalanskt: �ppet, Klassisk, 7.Ne5 Nc6 8.Nxc6
E05.9=Katalanskt: �ppet, Klassisk, 7.Qc2
E05.10=Katalanskt: �ppet, Klassisk Huvudvarianten
E05.11=Katalanskt: �ppet, Klassisk, 8.a4
E05.12=Katalanskt: �ppet, Klassisk, 8.a4 Bd7
E05.13=Katalanskt: �ppet, Klassisk, 8.a4 Bd7 9.Qxc4
E05.14=Katalanskt: �ppet, Klassisk, 8.a4 Bd7 9.Qxc4
E05.15=Katalanskt: �ppet, Klassisk, 8.a4, 10.Bg5 Bd5
E05.16=Katalanskt: �ppet, Klassisk, 8.a4, 10.Bg5 a5
E05.17=Katalanskt: �ppet, Klassisk, 8.Qxc4
E05.18=Katalanskt: �ppet, Klassisk, 8.Qxc4 b5 9.Qc2 Bb7
E05.19=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bg5
E05.20=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bd2
E05.21=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bd2 Be4
E05.22=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bf4
E05.23=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bf4 Nc6
E05.24=Katalanskt: �ppet, Klassisk, 8.Qxc4, 10.Bf4 Nc6 11.Rd1
E06.1=Katalanskt: St�ngt
E06.2=Katalanskt: St�ngt, 5.Nf3
E06.3=Katalanskt: St�ngt, 5.Nf3 O-O
E06.4=Katalanskt: St�ngt, 6.Qc2
E06.5=Katalanskt: St�ngt, 6.O-O
E06.6=Katalanskt: St�ngt, 6.O-O c5
E06.7=Katalanskt: St�ngt, 6.O-O c5 7.cxd5
E06.8=Katalanskt: St�ngt, 6.O-O c6
E06.9=Katalanskt: St�ngt, 6.O-O c6 7.b3
E06.10=Katalanskt: St�ngt, 6.O-O c6 7.Nbd2
E06.11=Katalanskt: St�ngt, 6.O-O c6 7.Nc3
E06.12=Katalanskt: St�ngt, 6.O-O c6 7.Nc3 b6
E06.13=Katalanskt: St�ngt, 6.O-O c6 7.Nc3 b6 8.Ne5
E06.14=Katalanskt: St�ngt, 6.O-O c6 7.Qc2
E06.15=Katalanskt: St�ngt, 6.O-O c6 7.Qc2 b6
E07.1=Katalanskt: St�ngt, 6...Nbd7
E07.2=Katalanskt: St�ngt, 6...Nbd7 7.Nbd2
E07.3=Katalanskt: St�ngt, 6...Nbd7 7.Qd3
E07.4=Katalanskt: St�ngt, 6...Nbd7 7.b3
E07.5=Katalanskt: St�ngt, 6...Nbd7 7.b3
E07.6=Katalanskt: St�ngt, 6...Nbd7 7.b3
E07.7=Katalanskt: St�ngt, 6...Nbd7 7.b3
E07.8=Katalanskt: St�ngt, 6...Nbd7 7.Nc3
E07.9=Katalanskt: St�ngt, 6...Nbd7 7.Nc3 dxc4
E07.10=Katalanskt: St�ngt, 6...Nbd7 7.Nc3 dxc4
E07.11=Katalanskt: St�ngt, 6...Nbd7 7.Nc3 c6
E07.12=Katalanskt: St�ngt, 6...Nbd7 7.Nc3 c6 8.Qb3
E07.13=Katalanskt: St�ngt, Botvinnikvarianten
E07.14=Katalanskt: St�ngt, 6...Nbd7 7.Nc3 c6 8.b3
E08.1=Katalanskt: St�ngt, 7.Qc2
E08.2=Katalanskt: St�ngt, 7.Qc2 c5
E08.3=Katalanskt: St�ngt, 7.Qc2 b6
E08.4=Katalanskt: St�ngt, 7.Qc2 c6
E08.5=Katalanskt: St�ngt, 7.Qc2 c6 8.Rd1
E08.6=Katalanskt: St�ngt, 7.Qc2 c6 8.Rd1 b6
E08.7=Katalanskt: St�ngt, Zagoryanskyvarianten
E08.8=Katalanskt: St�ngt, 7.Qc2 c6 8.Bf4
E08.9=Katalanskt: St�ngt, 7.Qc2 c6 8.Bf4 Nh5
E08.10=Katalanskt: St�ngt, 7.Qc2 c6 8.Bf4 Ne4
E08.11=Katalanskt: St�ngt, 7.Qc2 c6 8.Bf4 b6
E08.12=Katalanskt: St�ngt, 7.Qc2 c6 8.b3
E08.13=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b5
E08.14=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6
E08.15=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1
E08.16=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Ba6
E08.17=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Ba6 10.Nbd2
E08.18=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Bb7
E08.19=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Bb7 10.Nc3
E08.20=Katalanskt: St�ngt, Spasskys gambit
E08.21=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Bb7 10.Nc3 Rc8
E08.22=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Bb7 10.Nc3 Rc8 11.e4
E08.23=Katalanskt: St�ngt, 7.Qc2 c6 8.b3 b6 9.Rd1 Bb7 10.Nc3 Rc8 11.e4 dxe4
E09.1=Katalanskt: St�ngt, Huvudvarianten
E09.2=Katalanskt: St�ngt, Huvudvarianten, 8...b5
E09.3=Katalanskt: St�ngt, Huvudvarianten, 8...Re8
E09.4=Katalanskt: St�ngt, Huvudvarianten, 8...b6
E09.5=Katalanskt: St�ngt, Huvudvarianten, 9.b3
E09.6=Katalanskt: St�ngt, Huvudvarianten, Sokolskyvarianten
E09.7=Katalanskt: St�ngt, Huvudvarianten, 9.b3 Bb7
E09.8=Katalanskt: St�ngt, Huvudvarianten, 9.b3 Bb7 10.Bb2
E09.9=Katalanskt: St�ngt, Huvudvarianten, 9.b3 Bb7 10.Bb2 Rc8
E09.10=Katalanskt: St�ngt, Huvudvarianten, 9.e4
E09.11=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Ba6
E09.12=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Ba6 10.b3
E09.13=Katalanskt: St�ngt, Huvudvarianten, 9.e4 dxe4
E09.14=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Bb7
E09.15=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Bb7 10.e5
E09.16=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Bb7 10.b3
E09.17=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Bb7 10.b3 Rc8 11.Bb2
E09.18=Katalanskt: St�ngt, Huvudvarianten, 9.e4 Bb7 10.b3 Rc8 11.Bb2 c5
E10.1=Neoindiskt: 3.Nf3
E10.2=Neoindiskt: D�rys f�rsvar
E10.3=Neoindiskt: 3.Nf3 Be7
E10.4=Neoindiskt: 3.Nf3 a6
E10.5=Neoindiskt: 3.Nf3 a6 4.Nc3
E10.6=Neoindiskt: 3.Nf3 a6 4.Nc3 c5
E10.7=Neoindiskt: Blumenfeld/Benoni
E10.8=Neoindiskt: Blumenfeld/Benoni, 4.e3
E10.9=Neoindiskt: Blumenfeld/Benoni, 4.e3 b6
E10.10=Neoindiskt: Blumenfeld/Benoni, 4.e3 cxd4
E10.11=Blumenfelds motgambit
E10.12=Blumenfeld: 5.dxe6
E10.13=Blumenfeld: 5.dxe6 fxe6 6.cxb5
E10.14=Blumenfeld: 5.dxe6 fxe6 6.cxb5 d5
E10.15=Blumenfeld: 5.Bg5
E10.16=Blumenfeld: 5.Bg5 h6
E10.17=Blumenfeld: 5.Bg5 Qa5+
E10.18=Blumenfeld: 5.Bg5 exd5
E10.19=Blumenfeld: Spielmannvarianten
E11.1=Bogo-Indiskt
E11.2=Bogo-Indiskt: 4.Nbd2
E11.3=Bogo-Indiskt: 4.Nbd2 d5
E11.4=Bogo-Indiskt: 4.Nbd2 b6
E11.5=Bogo-Indiskt: 4.Nbd2 b6 5.a3
E11.6=Bogo-Indiskt: 4.Nbd2 b6 5.a3 Bxd2+
E11.7=Bogo-Indiskt: 4.Nbd2 b6 5.a3 Bxd2+ 6.Bxd2
E11.8=Bogo-Indiskt: 4.Nbd2 b6 5.a3 Bxd2+ 6.Bxd2 Bb7
E11.9=Bogo-Indiskt: 4.Nbd2 O-O
E11.10=Bogo-Indiskt: 4.Nbd2 O-O 5.a3
E11.11=Bogo-Indiskt: 4.Nbd2 O-O 5.a3 Bxd2+
E11.12=Bogo-Indiskt: 4.Nbd2 O-O 5.a3 Be7
E11.13=Bogo-Indiskt: Gr�nfeldvarianten
E11.14=Bogo-Indiskt: 4.Bd2
E11.15=Bogo-Indiskt: 4.Bd2 Be7
E11.16=Bogo-Indiskt: 4.Bd2 Be7 5.g3
E11.17=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5
E11.18=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2
E11.19=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2 O-O
E11.20=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2 O-O 7.O-O c6
E11.21=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2 O-O 7.O-O c6 8.Qc2
E11.22=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2 O-O 7.O-O c6 8.Qc2 b6
E11.23=Bogo-Indiskt: 4.Bd2 Be7 5.g3 d5 6.Bg2 O-O 7.O-O c6 8.Qc2 b6 9.Bf4
E11.24=Bogo-Indiskt: Vitolinvarianten
E11.25=Bogo-Indiskt: Vitolin, 6.g3
E11.26=Bogo-Indiskt: 4.Bd2 a5
E11.27=Bogo-Indiskt: 4.Bd2 a5 5.Nc3
E11.28=Bogo-Indiskt: 4.Bd2 a5 5.g3
E11.29=Bogo-Indiskt: Nimzowitschvarianten
E11.30=Bogo-Indiskt: Nimzowitsch, 5.Nc3
E11.31=Bogo-Indiskt: Nimzowitsch, 5.g3
E11.32=Bogo-Indiskt: Nimzowitsch, 5.g3 O-O
E11.33=Bogo-Indiskt: Nimzowitsch, 5.g3 O-O
E11.34=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6
E11.35=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Nc3
E11.36=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Nc3 Bxc3
E11.37=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Nc3 Bxc3 7.Bxc3
E11.38=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Nc3 Bxc3 7.Bxc3 Ne4
E11.39=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Nc3 Bxc3 7.Bxc3 Ne4 8.Rc1
E11.40=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Bg2
E11.41=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Bg2 Bxd2+
E11.42=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 6.Bg2 Bxd2+ 7.Nbxd2
E11.43=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 Huvudvarianten
E11.44=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 Huvudvarianten, 8...O-O
E11.45=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 Huvudvarianten, 8...a5
E11.46=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 Huvudvarianten, 8...a5 9.e4
E11.47=Bogo-Indiskt: Nimzowitsch, 5.g3 Nc6 Huvudvarianten, 8...a5 9.e4 e5 10.d5 Nb8
E11.48=Bogo-Indiskt: 4.Bd2 Bxd2+
E11.49=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Nbxd2
E11.50=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Qxd2
E11.51=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Qxd2 O-O
E11.52=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Qxd2 O-O 6.Nc3
E11.53=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Qxd2 O-O 6.Nc3 d5
E11.54=Bogo-Indiskt: 4.Bd2 Bxd2+ 5.Qxd2 O-O 6.Nc3 d5 7.e3
E12.1=Damindiskt
E12.2=Damindiskt: Milesvarianten
E12.3=Damindiskt: Miles, 5.e3 Be7
E12.4=Damindiskt: Miles, 5.e3 Be7 6.h3
E12.5=Damindiskt: Miles, 5.e3 Bb4+
E12.6=Damindiskt: Miles, 5.e3 Bb4+ 6.Nbd2
E12.7=Damindiskt: Miles, 5.e3 Bb4+ 6.Nfd2
E12.8=Damindiskt: Petrosian
E12.9=Damindiskt: Petrosian, 4...c5
E12.10=Damindiskt: Petrosian, 4...c5 5.d5
E12.11=Damindiskt: Petrosian, 4...c5 5.d5 Ba6
E12.12=Damindiskt: Petrosian, 4...c5 5.d5 Ba6 6.Qc2
E12.13=Damindiskt: Petrosian, 4...c5 5.d5 Ba6 6.Qc2 exd5 6.cxd5 g6
E12.14=Damindiskt: Petrosian, 4...Ba6
E12.15=Damindiskt: Petrosian, 4...Ba6 5.e3
E12.16=Damindiskt: Petrosian, 4...Ba6 5.Qc2
E12.17=Damindiskt: Petrosian, 4...Ba6 5.Qc2 c5
E12.18=Damindiskt: Petrosian, 4...Ba6 5.Qc2 Bb7
E12.19=Damindiskt: Petrosian, 4...Ba6 5.Qc2 Bb7 6.Nc3 c5
E12.20=Damindiskt: Petrosian, 4...Ba6 5.Qc2 Bb7 6.Nc3 c5 7.e4
E12.21=Damindiskt: Petrosian, 4...Ba6 5.Qc2 Bb7 6.Nc3 c5 7.e4 cd 8.Nxd4 Nc6
E12.22=Damindiskt: Petrosian, 4...Bb7
E12.23=Damindiskt: Petrosian, 5.Nc3
E12.24=Damindiskt: Petrosian, 5.Nc3 Bxf3
E12.25=Damindiskt: Petrosian, 5.Nc3 Be7
E12.26=Damindiskt: Petrosian, 5.Nc3 Ne4
E12.27=Damindiskt: Petrosian, 5.Nc3 g6
E12.28=Damindiskt: Petrosian, 5.Nc3 d5
E12.29=Damindiskt: Petrosian, 5.Nc3 d5 6.Bg5
E12.30=Damindiskt: Petrosian, 5.Nc3 d5 6.Bg5 Be7
E12.31=Damindiskt: Petrosian, 5.Nc3 d5 6.Bg5 Be7 7.Qa4+
E12.32=Damindiskt: Petrosian, 5.Nc3 d5 6.Bg5 Be7 7.Qa4+ c6
E12.33=Damindiskt: Petrosian, 5.Nc3 d5 6.Bg5 Be7 7.Qa4+ c6 8.Bxf6 Bxf6 9.cxd5 exd5
E12.34=Damindiskt: Petrosian, 6.cxd5 exd5
E12.35=Damindiskt: Petrosian, 6.cxd5 exd5 7.g3
E12.36=Damindiskt: Petrosian, 6.cxd5 exd5 7.Bg5
E12.37=Damindiskt: Petrosian, 6.cxd5 Nxd5
E12.38=Damindiskt: Petrosian, 6.cxd5 Nxd5 7.e4
E12.39=Damindiskt: Petrosian, 6.cxd5 Nxd5 7.e3
E12.40=Damindiskt: Petrosian, 6.cxd5 Nxd5 7.e3 g6
E12.41=Damindiskt: Petrosian, 6.cxd5 Nxd5 7.e3 Be7
E12.42=Damindiskt: Petrosian, Kasparov-varianten
E12.43=Damindiskt: Petrosian, Kasparov, 7...Be7
E12.44=Damindiskt: Petrosian, Kasparov, 7...c5
E12.45=Damindiskt: Petrosian, Kasparov, 7...Nxc3
E12.46=Damindiskt: Petrosian, Kasparov, 7...Nxc3 8.bxc3
E12.47=Damindiskt: Petrosian, Kasparov, 7...Nxc3 8.bxc3 c5
E12.48=Damindiskt: Petrosian, Kasparov, 7...Nxc3 8.bxc3 c5 9.e4
E12.49=Damindiskt: Petrosian, Kasparov, 7...Nxc3 8.bxc3 Be7
E12.50=Damindiskt: Petrosian, Kasparov, 7...Nxc3 8.bxc3 Be7 9.e4
E12.51=Damindiskt: 4.Bg5
E12.52=Damindiskt: 4.Nc3
E12.53=Damindiskt: 4.Nc3 Bb7
E12.54=Damindiskt: 4.Nc3 Bb7 5.Bg5
E12.55=Damindiskt: 5.Bg5 h6 6.Bh4 Be7
E12.56=Damindiskt: 5.Bg5 h6 6.Bh4 Be7 7.e3 Ne4
E12.57=Damindiskt: 5.Bg5 h6 6.Bh4 Be7 7.e3 c5
E12.58=Damindiskt: Botvinnikvarianten
E12.59=Damindiskt: Botvinnik, 8.Qc2
E12.60=Damindiskt: Botvinnik, 8.e3
E13.1=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4
E13.2=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.Qc2
E13.3=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.Qc2 g5
E13.4=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.Nd2
E13.5=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.Nd2 Bxc3
E13.6=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.Nd2 Bxc3 8.bxc3
E13.7=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3
E13.8=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 c5
E13.9=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+
E13.10=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3
E13.11=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3 d6
E13.12=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3 d6 9.Nd2
E13.13=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3 d6 9.Nd2 Nbd7
E13.14=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3 d6 9.Nd2 Nbd7 10.f3
E13.15=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 Bxc3+ 8.bxc3 d6 9.Nd2 Nbd7 10.f3 Qe7
E13.16=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5
E13.17=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5
E13.18=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4
E13.19=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2
E13.20=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2 Bxc3+
E13.21=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2 Bxc3+
E13.22=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2 Bxc3+ 10.bxc3 d6
E13.23=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2 Bxc3+ 10.bxc3 d6 11.Bd3
E13.24=Damindiskt: 5.Bg5 h6 6.Bh4 Bb4 7.e3 g5 8.Bg3 Ne4 9.Qc2 Bxc3+ 10.bxc3 d6 11.Bd3 f5
E14.1=Damindiskt: 4.e3
E14.2=Damindiskt: 4.e3 Bb4+
E14.3=Damindiskt: 4.e3 Bb7
E14.4=Damindiskt: 4.e3 Bb7 5.Nc3
E14.5=Damindiskt: 4.e3 Bb7 5.Nc3 d5
E14.6=Damindiskt: 4.e3 Bb7 5.Bd3
E14.7=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+
E14.8=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2
E14.9=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2 c5
E14.10=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2 O-O
E14.11=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2 O-O 7.O-O d5
E14.12=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2 O-O 7.O-O d5 8.a3
E14.13=Damindiskt: 4.e3 Bb7 5.Bd3 Bb4+ 6.Nbd2 O-O 7.O-O d5 8.a3 Be7
E14.14=Damindiskt: Dreevvarianten
E14.15=Damindiskt: 4.e3 Bb7 5.Bd3 Be7
E14.16=Damindiskt: 4.e3 Bb7 5.Bd3 Be7 6.O-O
E14.17=Damindiskt: 4.e3 Bb7 5.Bd3 Be7 6.O-O O-O
E14.18=Damindiskt: 4.e3 Bb7 5.Bd3 Be7 6.O-O O-O 7.Nc3
E14.19=Damindiskt: 4.e3 Bb7 5.Bd3 d5
E14.20=Damindiskt: 4.e3 Bb7 5.Bd3 d5 6.O-O
E14.21=Damindiskt: 4.e3 Bb7 5.Bd3 d5 6.O-O Bd6
E14.22=Damindiskt: 4.e3 Bb7 5.Bd3 d5 6.O-O Bd6 7.b3
E14.23=Damindiskt: 4.e3 Bb7 5.Bd3 d5 6.O-O Bd6 7.Nc3
E14.24=Damindiskt: 4.e3 Bb7 5.Bd3 c5
E14.25=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.Nc3
E14.26=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O
E14.27=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O cxd4
E14.28=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O cxd4 7.exd4
E14.29=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7
E14.30=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nbd2
E14.31=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3
E14.32=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3
E14.33=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3 O-O 8.Bb2 d5
E14.34=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3 O-O 8.Bb2 cxd4
E14.35=Damindiskt: Averbakhvarianten
E14.36=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3 O-O 8.Bb2 cxd4 9.exd4
E14.37=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.b3 O-O 8.Bb2 cxd4 9.exd4 d5
E14.38=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nc3
E14.39=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nc3 O-O
E14.40=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nc3 cxd4
E14.41=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nc3 cxd4 8.exd4
E14.42=Damindiskt: 4.e3 Bb7 5.Bd3 c5 6.O-O Be7 7.Nc3 cxd4 8.exd4 d5
E15.1=Damindiskt: 4.g3
E15.2=Damindiskt: 4.g3 Bb4+
E15.3=Damindiskt: 4.g3 Bb4+
E15.4=Damindiskt: 4.g3 Bb4+ 5.Bd2 Bxd2+
E15.5=Damindiskt: 4.g3 Bb4+ 5.Bd2 Bxd2+ 6.Qxd2 Ba6
E15.6=Damindiskt: Nimzowitschvarianten (4.g3 Ba6)
E15.7=Damindiskt: Nimzowitsch, 5.Qb3
E15.8=Damindiskt: Nimzowitsch, 5.Qc2
E15.9=Damindiskt: Nimzowitsch, 5.Nbd2
E15.10=Damindiskt: Nimzowitsch, 5.Nbd2 c5
E15.11=Damindiskt: Nimzowitsch, 5.Nbd2 Bb7
E15.12=Damindiskt: Nimzowitsch, 5.Nbd2 Bb7 6.Bg2
E15.13=Damindiskt: Nimzowitsch, 5.Nbd2 Bb7 6.Bg2 c5
E15.14=Damindiskt: Nimzowitsch, 5.Nbd2 Bb4
E15.15=Damindiskt: Nimzowitsch, 5.Qa4
E15.16=Damindiskt: Nimzowitsch, 5.Qa4 Be7
E15.17=Damindiskt: Nimzowitsch, 5.Qa4 c6
E15.18=Damindiskt: Nimzowitsch, 5.Qa4 c6 6.Nc3 b5
E15.19=Damindiskt: Nimzowitsch, 5.Qa4 c5
E15.20=Damindiskt: Nimzowitsch, 5.Qa4 c5 6.Bg2 Bb7
E15.21=Damindiskt: Nimzowitsch, 5.Qa4 c5 6.Bg2 Bb7 7.dxc5
E15.22=Damindiskt: Nimzowitsch, 5.Qa4 c5 6.Bg2 Bb7 7.O-O
E15.23=Damindiskt: Nimzowitsch, 5.b3 
E15.24=Damindiskt: Nimzowitsch, 5.b3 b5
E15.25=Damindiskt: Nimzowitsch, 5.b3 b5 6.cxb5
E15.26=Damindiskt: Nimzowitsch, 5.b3 d5
E15.27=Damindiskt: Nimzowitsch, 5.b3 d5 6.cxd5
E15.28=Damindiskt: Nimzowitsch, 5.b3 d5 6.Bg2
E15.29=Damindiskt: Nimzowitsch, 5.b3 Bb7
E15.30=Damindiskt: Nimzowitsch, 5.b3 Bb7 6.Bg2
E15.31=Damindiskt: Nimzowitsch, 5.b3 Bb7, 7...a5
E15.32=Damindiskt: Nimzowitsch, 5.b3 Bb7, 7...a5 8.O-O O-O
E15.33=Damindiskt: Nimzowitsch, 5.b3 Bb4+
E15.34=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7
E15.35=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Nc3
E15.36=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2
E15.37=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2 d5
E15.38=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2 d5
E15.39=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2 c6
E15.40=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2 c6 8.O-O
E15.41=Damindiskt: Nimzowitsch, 5.b3 Bb4+ 6.Bd2 Be7 7.Bg2 c6 8.O-O d5
E15.42=Damindiskt: Nimzowitsch, 5.b3 Bb4+, Huvudvarianten
E15.43=Damindiskt: Nimzowitsch, 5.b3 Bb4+, Huvudvarianten, 9.Ne5
E15.44=Damindiskt: Nimzowitsch, 5.b3 Bb4+, Huvudvarianten, 9.Ne5 Nfd7
E15.45=Damindiskt: 4.g3 Bb7
E15.46=Damindiskt: 4.g3 Bb7
E15.47=Damindiskt: 4.g3 Bb7 5.Bg2 Qc8
E15.48=Damindiskt: 4.g3 Bb7 5.Bg2 Qc8 6.O-O c5 7.d5
E15.49=Damindiskt: 4.g3 Bb7 5.Bg2 c5
E15.50=Damindiskt: Buergervarianten
E15.51=Damindiskt: Rubinsteinvarianten
E16.1=Damindiskt: Capablancavarianten
E16.2=Damindiskt: Capablanca, 6.Nbd2
E16.3=Damindiskt: Capablanca, 6.Nbd2 O-O
E16.4=Damindiskt: Capablanca, 6.Nbd2 O-O 7.O-O d5
E16.5=Damindiskt: Capablanca, 6.Bd2
E16.6=Damindiskt: Capablanca, 6.Bd2 c5
E16.7=Damindiskt: Capablanca, Yates-varianten
E16.8=Damindiskt: Capablanca, Yates, 7.O-O O-O
E16.9=Damindiskt: Capablanca, Nimzowitsch-varianten
E16.10=Damindiskt: Capablanca, Nimzowitsch, 7.O-O Bxd2 8.Qxd2
E16.11=Damindiskt: Capablanca, Riumin-varianten
E16.12=Damindiskt: Capablanca, Riumin, 7.Nc3
E16.13=Damindiskt: Capablanca, Riumin, 7.Nc3 O-O
E16.14=Damindiskt: Capablanca, Riumin, 7.Nc3 O-O 8.O-O
E16.15=Damindiskt: Capablanca, Riumin, 7.Nc3 O-O 8.O-O d5
E16.16=Damindiskt: Capablanca, 6...Bxd2+
E16.17=Damindiskt: Capablanca, 6...Bxd2+ 7.Nbxd2
E16.18=Damindiskt: Capablanca, 6...Bxd2+ 7.Qxd2
E16.19=Damindiskt: Capablanca, 6...Bxd2+ 7.Qxd2 O-O
E16.20=Damindiskt: Capablanca, 6...Bxd2+ 7.Qxd2 O-O 8.O-O
E16.21=Damindiskt: Capablanca, 6...Bxd2+ 7.Qxd2 O-O 8.Nc3
E17.1=Damindiskt: 5.Bg2 Be7
E17.2=Damindiskt: 6.Nc3
E17.3=Damindiskt: 6.Nc3 d5
E17.4=Damindiskt: 6.Nc3 O-O
E17.5=Damindiskt: 6.Nc3 O-O 7.Qc2
E17.6=Damindiskt: 6.Nc3 O-O 7.Qc2 c5
E17.7=Damindiskt: 6.Nc3 O-O 7.Qc2 d5
E17.8=Damindiskt: 6.Nc3 Ne4
E17.9=Damindiskt: 6.Nc3 Ne4 7.Qc2
E17.10=Damindiskt: Opovcenskyvarianten
E17.11=Damindiskt: Opovcensky, 7...O-O
E17.12=Damindiskt: Opovcensky, 7...f5
E17.13=Damindiskt: Opovcensky, 7...Bf6
E17.14=Damindiskt: 6.O-O
E17.15=Damindiskt: 6.O-O d5
E17.16=Damindiskt: 6.O-O O-O
E17.17=Damindiskt: 6.O-O O-O 7.Qc2
E17.18=Damindiskt: 6.O-O O-O 7.Re1
E17.19=Damindiskt: 6.O-O O-O 7.Re1 d5
E17.20=Damindiskt: Euwevarianten
E17.21=Damindiskt: Euwe, 7...c5
E17.22=Damindiskt: Euwe, 7...d5
E17.23=Damindiskt: Pomarvarianten
E17.24=Damindiskt: Pomar, 7...exd5
E17.25=Damindiskt: Pomar, Taimanovvarianten
E17.26=Damindiskt: Pomar, Polugaevskyvarianten
E17.27=Damindiskt: Pomar, Polugaevsky, 8...c6
E17.28=Damindiskt: Pomar, Polugaevsky, 8...c6 9.cxd5 Nxd5
E17.29=Damindiskt: Pomar, Polugaevsky, 8...c6 9.cxd5 Nxd5 10.Nf5 Nc7
E17.30=Damindiskt: Pomar, Polugaevsky, 8...c6 9.cxd5 Nxd5 10.Nf5 Nc7 11.e4
E18.1=Damindiskt: 7.Nc3
E18.2=Damindiskt: 7.Nc3 c5
E18.3=Damindiskt: 7.Nc3 d6
E18.4=Damindiskt: 7.Nc3 Na6
E18.5=Damindiskt: 7.Nc3 d5
E18.6=Damindiskt: 7.Nc3 d5 8.cxd5
E18.7=Damindiskt: 7.Nc3 d5 8.cxd5 exd5
E18.8=Damindiskt: 7.Nc3 d5 8.Ne5
E18.9=Damindiskt: 7.Nc3 d5 8.Ne5 c6
E18.10=Damindiskt: 7.Nc3 d5 8.Ne5 Nbd7
E18.11=Damindiskt: 7.Nc3 d5 8.Ne5 Na6
E18.12=Damindiskt: 7.Nc3 d5 8.Ne5 Na6 9.cxd5 exd5
E18.13=Damindiskt: 7.Nc3 Ne4
E18.14=Damindiskt: 7.Nc3 Ne4 8.Bd2
E18.15=Damindiskt: 7.Nc3 Ne4 8.Bd2 d5
E18.16=Damindiskt: 7.Nc3 Ne4 8.Bd2 d5 9.cxd5 exd5
E18.17=Damindiskt: 7.Nc3 Ne4 8.Bd2 f5
E18.18=Damindiskt: 7.Nc3 Ne4 8.Bd2 f5 9.d5
E18.19=Damindiskt: 7.Nc3 Ne4 8.Bd2 f5 9.d5 Bf6
E18.20=Damindiskt: 7.Nc3 Ne4 8.Bd2 f5 9.d5 Bf6 10.Rc1
E18.21=Damindiskt: 7.Nc3 Ne4 8.Bd2 Bf6
E18.22=Damindiskt: 7.Nc3 Ne4 8.Bd2 Bf6 9.Rc1
E18.23=Damindiskt: 7.Nc3 Ne4 8.Nxe4
E18.24=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.d5
E18.25=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Bf4
E18.26=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Nh4
E18.27=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1
E18.28=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1 Bxg2 10.Nxg2
E18.29=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1 Bxg2 10.Nxg2 d5
E18.30=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1 Bxg2 10.Nxg2 d5 11.Qa4
E18.31=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1 Bxg2 10.Nxg2 d5 11.Qa4 Qd7
E18.32=Damindiskt: 7.Nc3 Ne4 8.Nxe4 Bxe4 9.Ne1 Bxg2 10.Nxg2 d5 11.Qa4 dxc4
E18.33=Damindiskt: Gamla huvudvarianten, 8.Qc2
E18.34=Damindiskt: Gamla huvudvarianten, 8.Qc2 Nxc3
E18.35=Damindiskt: Gamla huvudvarianten, 8.Qc2 Nxc3 9.bxc3
E19.1=Damindiskt: Gamla huvudvarianten, 9.Qxc3
E19.2=Damindiskt: Gamla huvudvarianten, 9.Qxc3 d6
E19.3=Damindiskt: Gamla huvudvarianten, 9.Qxc3 d6 10.b3
E19.4=Damindiskt: Gamla huvudvarianten, 9.Qxc3 Be4
E19.5=Damindiskt: Gamla huvudvarianten, 9.Qxc3 Be4 10.Ne1
E19.6=Damindiskt: Gamla huvudvarianten, 9.Qxc3 f5
E19.7=Damindiskt: Gamla huvudvarianten, 9.Qxc3 f5 10.Rd1
E19.8=Damindiskt: Gamla huvudvarianten, 9.Qxc3 f5 10.b3
E19.9=Damindiskt: Gamla huvudvarianten, 9.Qxc3 f5 10.b3 Bf6 11.Bb2 d6
E19.10=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5
E19.11=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.b3
E19.12=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1
E19.13=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1 d6
E19.14=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1 d6 11.b3
E19.15=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1 d6 11.b3 Bf6
E19.16=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1 d6 11.b3 Bf6
E19.17=Damindiskt: Gamla huvudvarianten, 9.Qxc3 c5 10.Rd1 d6 11.b3 Bf6 12.Bb2 Qe7
E20.1=Nimzoindiskt f�rsvar
E20.2=Nimzoindiskt: Mikenas attack
E20.3=Nimzoindiskt: 4.Bd2
E20.4=Nimzoindiskt: 4.Bd2 O-O
E20.5=Nimzoindiskt: 4.Bd2 O-O 5.Nf3
E20.6=Nimzoindiskt: Romanishin
E20.7=Nimzoindiskt: Romanishin, 4...c5
E20.8=Nimzoindiskt: Romanishin, 4...c5 5.d5
E20.9=Nimzoindiskt: Romanishin, 4...c5 5.Nf3
E20.10=Nimzoindiskt: Romanishin, 4...c5 5.Nf3 Ne4
E20.11=Nimzoindiskt: Romanishin, 4...c5 5.Nf3 Nc6
E20.12=Nimzoindiskt: Romanishin, 4...c5 5.Nf3 O-O
E20.13=Nimzoindiskt: Romanishin, 4...c5 5.Nf3 cxd4
E20.14=Nimzoindiskt: Romanishin, 6.Nxd4
E20.15=Nimzoindiskt: Romanishin, 6.Nxd4 O-O
E20.16=Nimzoindiskt: Romanishin, 6.Nxd4 O-O 7.Bg2
E20.17=Nimzoindiskt: Romanishin, 6.Nxd4 O-O 7.Bg2 d5
E20.18=Nimzoindiskt: Romanishin, 8.cxd5
E20.19=Nimzoindiskt: 4.f3 (Kmoch)
E20.20=Nimzoindiskt: 4.f3 d5
E20.21=Nimzoindiskt: 4.f3 d5 5.a3 Be7
E20.22=Nimzoindiskt: 4.f3 c5
E20.23=Nimzoindiskt: 4.f3 c5 5.d5
E21.1=Nimzoindiskt: Tre springare
E21.2=Nimzoindiskt: Nimzo-damhybrid
E21.3=Nimzoindiskt: Nimzo-damhybrid, 5.Qc2
E21.4=Nimzoindiskt: Nimzo-damhybrid, 5.Qc2 Bb7
E21.5=Nimzoindiskt: Nimzo-damhybrid, 5.Qb3
E21.6=Nimzoindiskt: Nimzo-damhybrid, 5.Qb3 a5
E21.7=Nimzoindiskt: Nimzo-damhybrid, 5.Qb3 c5
E21.8=Nimzoindiskt: Nimzo-damhybrid, 5.Bg5
E21.9=Nimzoindiskt: Nimzo-damhybrid, 5.Bg5 Bb7
E21.10=Nimzoindiskt: Tre springare, 4...O-O
E21.11=Nimzoindiskt: Tre springare, 4...Bxc3+
E21.12=Nimzoindiskt: Tre springare, 4...c5
E21.13=Nimzoindiskt: Tre springare, Euwevarianten
E22.1=Nimzoindiskt: Spielmannvarianten
E22.2=Nimzoindiskt: Spielmann, 4...Nc6
E22.3=Nimzoindiskt: Spielmann, 4...c5
E22.4=Nimzoindiskt: Spielmann, 4...c5 5.Nf3
E22.5=Nimzoindiskt: Spielmann, 4...c5 5.dxc5
E22.6=Nimzoindiskt: Spielmann, 4...c5 5.dxc5 Na6
E23.1=Nimzoindiskt: Spielmann, 4...c5 5.dxc5 Nc6
E23.3=Nimzoindiskt: Spielmann, San Removarianten
E23.4=Nimzoindiskt: Spielmann, St�hlbergvarianten
E23.2=Nimzoindiskt: Spielmann, Carlsbadvarianten
E24.1=Nimzoindiskt: S�misch
E24.2=Nimzoindiskt: S�misch
E24.3=Nimzoindiskt: S�misch, 5...b6
E24.4=Nimzoindiskt: S�misch, 5...b6 6.f3
E24.5=Nimzoindiskt: S�misch, 5...d5
E24.6=Nimzoindiskt: S�misch, 5...d5 6.f3
E24.7=Nimzoindiskt: S�misch, 5...c5
E24.8=Nimzoindiskt: S�misch, 5...c5 6.f3
E24.9=Nimzoindiskt: S�misch, 5...c5 6.f3 d5
E24.10=Nimzoindiskt: S�misch, Botvinnikvarianten
E25.1=Nimzoindiskt: S�misch, 5...c5 6.f3 d5 7.cxd5
E25.2=Nimzoindiskt: S�misch, 5...c5 6.f3 d5 7.cxd5 Nxd5
E25.3=Nimzoindiskt: S�misch, 5...c5 6.f3 d5 7.cxd5 Nxd5 8.Qd3
E25.4=Nimzoindiskt: S�misch, Keresvarianten
E25.5=Nimzoindiskt: S�misch, Keres, Romanovskyvarianten
E25.6=Nimzoindiskt: S�misch, Keres, Romanovsky, 9.e4
E25.7=Nimzoindiskt: S�misch, Keres, Romanovsky, 9.Nh3
E26.1=Nimzoindiskt: S�misch, 5...c5 6.e3
E26.3=Nimzoindiskt: S�misch, O'Kellyvarianten
E26.2=Nimzoindiskt: S�misch, 5...c5 6.e3 Nc6
E27.1=Nimzoindiskt: S�misch, 5...O-O
E27.2=Nimzoindiskt: S�misch, 5...O-O 6.f3
E27.3=Nimzoindiskt: S�misch, 5...O-O 6.f3 d5
E28.1=Nimzoindiskt: S�misch, 5...O-O 6.e3
E28.2=Nimzoindiskt: S�misch, 5...O-O 6.e3
E28.3=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5
E28.4=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Ne2
E28.5=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Bd3
E28.6=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Bd3 b6
E29.1=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Bd3 Nc6
E29.2=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Bd3 Nc6 8.Ne2
E29.3=Nimzoindiskt: S�misch, 5...O-O 6.e3 c5 7.Bd3 Nc6 8.Ne2 b6
E29.4=Nimzoindiskt: S�misch, Capablancavarianten
E30.1=Nimzoindiskt: Leningrad
E30.2=Nimzoindiskt: Leningrad, 4...O-O
E30.3=Nimzoindiskt: Leningrad, 4...c5
E30.4=Nimzoindiskt: Leningrad, 4...c5 5.d5
E30.5=Nimzoindiskt: Leningrad, 4...c5 5.d5 exd5
E30.6=Nimzoindiskt: Leningrad, 4...c5 5.d5 Bxc3+
E30.7=Nimzoindiskt: Leningrad, 4...c5 5.d5 d6
E30.8=Nimzoindiskt: Leningrad, 4...c5 5.d5 d6 6.e3
E30.9=Nimzoindiskt: Leningrad, 4...c5 5.d5 h6
E30.10=Nimzoindiskt: Leningrad, 4...h6
E30.11=Nimzoindiskt: Leningrad, 4...h6 5.Bxf6
E30.12=Nimzoindiskt: Leningrad, 4...h6 5.Bh4
E30.13=Nimzoindiskt: Leningrad, 4...h6 5.Bh4 c5
E30.14=Nimzoindiskt: Leningrad, 6.d5
E30.15=Nimzoindiskt: Leningrad, 6.d5 exd5
E30.16=Nimzoindiskt: Leningrad, 6.d5 exd5
E30.17=Nimzoindiskt: Leningrad, 6.d5 b5 gambit
E30.18=Nimzoindiskt: Leningrad, 6.d5 Bxc3+
E31.1=Nimzoindiskt: Leningrad, Huvudvarianten
E31.2=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3
E31.3=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 g5
E31.4=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 exd5
E31.5=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 e5
E31.7=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 Qe7
E31.6=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 O-O
E31.8=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 Bxc3+
E31.9=Nimzoindiskt: Leningrad, Huvudvarianten, 7.e3 Bxc3+
E31.10=Nimzoindiskt: Leningrad, Huvudvarianten, 8...Qe7
E31.11=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5
E31.12=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5 9.Nf3
E31.13=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5 9.Qc2
E31.14=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5 9.Bd3
E31.15=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5 9.f3
E31.16=Nimzoindiskt: Leningrad, Huvudvarianten, 8...e5 9.f3 Nbd7
E32.1=Nimzoindiskt: Klassiska varianten
E32.2=Nimzoindiskt: Klassisk, 4...b6
E32.3=Nimzoindiskt: Klassisk, 4...d6
E32.4=Nimzoindiskt: Klassisk, 4...O-O
E32.5=Nimzoindiskt: Klassisk, 4...O-O 5.Bg5
E32.6=Nimzoindiskt: Klassisk, 4...O-O 5.e4
E32.7=Nimzoindiskt: Klassisk, 4...O-O 5.Nf3
E32.8=Nimzoindiskt: Klassisk, 4...O-O 5.a3
E32.9=Nimzoindiskt: Klassisk, 4...O-O 5.a3
E32.10=Nimzoindiskt: Klassisk, 4...O-O 5.a3
E32.11=Nimzoindiskt: Klassisk, Adorjans gambit
E32.12=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...d6
E32.13=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...Ne4
E32.14=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6
E32.15=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Nf3
E32.16=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5
E32.17=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Ba6
E32.18=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7
E32.19=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7 8.f3
E32.20=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7 8.f3 h6
E32.21=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7 8.f3 h6 9.Bh4
E32.22=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7 8.e3
E32.23=Nimzoindiskt: Klassisk, 4...O-O 5.a3, 6...b6 7.Bg5 Bb7 8.e3 d6
E33.1=Nimzoindiskt: Klassisk, 4...Nc6
E33.2=Nimzoindiskt: Klassisk, 4...Nc6 5.Nf3
E33.3=Nimzoindiskt: Klassisk, 4...Nc6 5.Nf3 d5
E33.4=Nimzoindiskt: Klassisk, Milner-Barry (Zurich)varianten
E33.5=Nimzoindiskt: Klassisk, Milner-Barry (Zurich), 6.a3
E33.6=Nimzoindiskt: Klassisk, Milner-Barry (Zurich), 6.a3 Bxc3+ 7.Qxc3
E33.7=Nimzoindiskt: Klassisk, Milner-Barry (Zurich), 6.Bd2
E33.8=Nimzoindiskt: Klassisk, Milner-Barry (Zurich), 6.Bd2 O-O
E34.1=Nimzoindiskt: Klassisk, Noavarianten
E34.2=Nimzoindiskt: Klassisk, Noa, 5.e3
E34.3=Nimzoindiskt: Klassisk, Noa, 5.e3 O-O
E34.4=Nimzoindiskt: Klassisk, Noa, 5.cxd5
E34.5=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5
E34.6=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.e3
E34.7=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.e3 c5
E34.8=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.Nf3
E34.9=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.Nf3 c5
E34.10=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.Nf3 Qf5
E34.11=Nimzoindiskt: Klassisk, Noa, 5.cxd5 Qxd5 6.Nf3 Qf5 7.Qb3
E34.12=Nimzoindiskt: Klassisk, Noa, Dambyte
E35.1=Nimzoindiskt: Klassisk, Noa, Avbyte
E35.2=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.a3
E35.3=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5
E35.4=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5 c5
E35.5=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5 h6
E35.6=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5 h6 7.Bh4
E35.7=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5 h6 7.Bh4 c5
E35.8=Nimzoindiskt: Klassisk, Noa, Avbyte, 6.Bg5 h6 7.Bxf6
E36.1=Nimzoindiskt: Klassisk, Noa, 5.a3
E36.2=Nimzoindiskt: Klassisk, Noa, 5.a3 Be7
E36.3=Nimzoindiskt: Klassisk, Noa, 5.a3 Bxc3+
E36.4=Nimzoindiskt: Klassisk, Noa, 5.a3 Bxc3+
E36.5=Nimzoindiskt: Klassisk, Noa, 5.a3 Bxc3+ 6.Qxc3 dxc4
E36.6=Nimzoindiskt: Klassisk, Noa, 5.a3 Bxc3+ 6.Qxc3 O-O
E36.7=Nimzoindiskt: Klassisk, Noa, Botvinnikvarianten
E36.8=Nimzoindiskt: Klassisk, Noa, Huvudvarianten
E37.1=Nimzoindiskt: Klassisk, Noa, Huvudvarianten, 7.Qc2
E37.2=Nimzoindiskt: Klassisk, Noa, Huvudvarianten, 7.Qc2 Nc6
E37.3=Nimzoindiskt: Klassisk, Noa, San Removarianten
E37.4=Nimzoindiskt: Klassisk, Noa, Huvudvarianten, 7.Qc2 c5
E37.5=Nimzoindiskt: Klassisk, Noa, Huvudvarianten, 7.Qc2 c5 8.dxc5 Nc6
E38.1=Nimzoindiskt: Klassisk, 4...c5
E38.2=Nimzoindiskt: Klassisk, 4...c5 5.Nf3
E38.3=Nimzoindiskt: Klassisk, 4...c5 5.e3
E38.4=Nimzoindiskt: Klassisk, 4...c5 5.dxc5
E38.5=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Bxc5
E38.6=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Bxc5 6.Nf3
E38.7=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Bxc5 6.Nf3 Qb6
E38.8=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Qc7
E38.9=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Nc6
E38.10=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6
E38.11=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6 6.a3 Bxc3+ 7.Qxc3
E38.12=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6: 8.b4
E38.13=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6: 8.b4 Nce4
E38.14=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6: 8.b4 Nce4 9.Qd4
E38.15=Nimzoindiskt: Klassisk, 4...c5 5.dxc5 Na6: 8.b4 Nce4 9.Qd4 d5 10.c5
E39.1=Nimzoindiskt: Klassisk, Pircvarianten
E39.2=Nimzoindiskt: Klassisk, Pirc, 6.Bf4
E39.3=Nimzoindiskt: Klassisk, Pirc, 6.Nf3
E39.4=Nimzoindiskt: Klassisk, Pirc, 6.Nf3 Bxc5
E39.5=Nimzoindiskt: Klassisk, Pirc, 6.Nf3 Na6
E39.6=Nimzoindiskt: Klassisk, Pirc, 6.Nf3 Na6 7.Bd2
E39.7=Nimzoindiskt: Klassisk, Pirc, 6.Nf3 Na6 7.a3
E39.8=Nimzoindiskt: Klassisk, Pirc, 6.Nf3 Na6 7.g3
E39.9=Nimzoindiskt: Klassisk, Pirc, 6.a3
E39.10=Nimzoindiskt: Klassisk, Pirc, 6.a3 Bxc5 7.Nf3
E39.11=Nimzoindiskt: Klassisk, Pirc, 6.a3 Bxc5 7.Nf3 Nc6
E39.12=Nimzoindiskt: Klassisk, Pirc, 6.a3 Bxc5 7.Nf3 b6
E39.13=Nimzoindiskt: Klassisk, Pirc, 6.a3 Bxc5 7.Nf3 b6 8.Bg5
E40.1=Nimzoindiskt: Rubinstein
E40.2=Nimzoindiskt: Taimanov
E40.3=Nimzoindiskt: Taimanov, 5.Ne2
E40.4=Nimzoindiskt: Taimanov, 5.Ne2 d5
E40.5=Nimzoindiskt: Taimanov, 5.Bd3
E41.1=Nimzoindiskt: 4.e3 c5
E41.2=Nimzoindiskt: 4.e3 c5 5.Nf3
E41.3=Nimzoindiskt: 4.e3 c5 5.Bd3
E41.4=Nimzoindiskt: 4.e3 c5 5.Bd3 Nc6
E41.5=Nimzoindiskt: 4.e3 c5 5.Bd3 Nc6 6.Ne2
E41.6=Nimzoindiskt: 4.e3 c5 5.Bd3 Nc6 6.Nf3
E41.7=Nimzoindiskt: 4.e3 c5, H�bnervarianten
E41.8=Nimzoindiskt: H�bner, 8.e4
E41.9=Nimzoindiskt: H�bner, 8.e4 e5 9.d5 Ne7
E41.10=Nimzoindiskt: H�bner, 8.O-O
E41.11=Nimzoindiskt: H�bner, 8.O-O e5
E41.12=Nimzoindiskt: H�bner, 8.O-O e5 9.Nd2
E42.1=Nimzoindiskt: 4.e3 c5 5.Ne2
E42.2=Nimzoindiskt: 4.e3 c5 5.Ne2 d5
E42.3=Nimzoindiskt: 4.e3 c5 5.Ne2 cxd4 6.exd4
E42.4=Nimzoindiskt: 4.e3 c5 5.Ne2 cxd4 6.exd4 d5
E42.5=Nimzoindiskt: 4.e3 c5 5.Ne2 cxd4 6.exd4 O-O
E42.6=Nimzoindiskt: 4.e3 c5 5.Ne2 cxd4 6.exd4 O-O 7.a3 Be7
E43.1=Nimzoindiskt: Nimzowitsch (Fischer)varianten
E43.2=Nimzoindiskt: Nimzowitsch, 5.Bd3
E43.3=Nimzoindiskt: Nimzowitsch, 5.Nf3
E43.4=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7
E43.5=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7 6.Bd3
E43.6=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7 6.Bd3 O-O
E43.7=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7 6.Bd3 O-O 7.O-O
E43.8=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7 6.Bd3 Ne4
E43.9=Nimzoindiskt: Nimzowitsch, 5.Nf3 Bb7 6.Bd3 Ne4 7.O-O
E43.10=Nimzoindiskt: Nimzowitsch, Keene-varianten
E44.1=Nimzoindiskt: Nimzowitsch, 5.Ne2
E44.2=Nimzoindiskt: Nimzowitsch, 5.Ne2 Bb7
E44.3=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ne4
E44.4=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ne4 6.Bd2
E44.5=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ne4 6.Qc2
E45.1=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6
E45.2=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.a3
E45.3=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.a3 Be7
E45.4=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.a3 Bxc3+
E45.5=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.Ng3
E45.6=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.Ng3 h5
E45.7=Nimzoindiskt: Nimzowitsch, 5.Ne2 Ba6 6.Ng3 Bxc3+
E46.1=Nimzoindiskt: 4.e3 O-O
E46.2=Nimzoindiskt: Reshevskyvarianten
E46.3=Nimzoindiskt: Reshevskyvarianten
E46.4=Nimzoindiskt: Reshevskyvarianten
E46.5=Nimzoindiskt: Reshevskyvarianten
E46.6=Nimzoindiskt: Reshevsky, Simagin-varianten
E46.7=Nimzoindiskt: Reshevsky, 6.a3 Be7
E46.8=Nimzoindiskt: Reshevsky, 6.a3 Be7 7.cxd5
E46.9=Nimzoindiskt: Reshevsky, 6.a3 Be7 7.cxd5 exd5
E47.1=Nimzoindiskt: 4.e3 O-O 5.Bd3
E47.2=Nimzoindiskt: 4.e3 O-O 5.Bd3 b6
E47.3=Nimzoindiskt: 4.e3 O-O 5.Bd3 d6
E47.4=Nimzoindiskt: 4.e3 O-O 5.Bd3 c5
E47.5=Nimzoindiskt: 4.e3 O-O 5.Bd3 c5 6.Ne2
E47.6=Nimzoindiskt: 4.e3 O-O 5.Bd3 c5 6.Ne2 cxd4
E48.1=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5
E48.2=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.cxd5
E48.3=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2
E48.4=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5
E48.5=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.O-O
E48.6=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.O-O cxd4 8.exd4
E48.7=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.cxd5
E48.8=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.cxd5 cxd4 8.exd4
E48.9=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.cxd5 cxd4 8.exd4 Nxd5
E48.10=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.Ne2 c5 7.cxd5 cxd4 8.exd4 Nxd5 9.O-O
E48.11=Nimzoindiskt: 4.e3 O-O 5.Bd3 d5 6.a3
E49.1=Nimzoindiskt: Botvinniks system
E49.2=Nimzoindiskt: Botvinnik, 7...dxc4
E49.3=Nimzoindiskt: Botvinnik, 7...dxc4 8.Bxc4 c5
E49.4=Nimzoindiskt: Botvinnik, 7...dxc4 8.Bxc4 c5 9.Ne2
E49.5=Nimzoindiskt: Botvinnik, 7...c5
E49.6=Nimzoindiskt: Botvinnik, 7...c5 8.cxd5
E49.7=Nimzoindiskt: Botvinnik, 7...c5 8.cxd5 exd5 9.Ne2
E49.8=Nimzoindiskt: Botvinnik, 7...c5 8.cxd5 exd5
E50.1=Nimzoindiskt: 4.e3 O-O 5.Nf3
E50.2=Nimzoindiskt: 4.e3 O-O 5.Nf3 Ne4
E50.3=Nimzoindiskt: 4.e3 O-O 5.Nf3 b6
E50.4=Nimzoindiskt: 4.e3 O-O 5.Nf3 c5
E50.5=Nimzoindiskt: 4.e3 O-O 5.Nf3 c5 6.Bd3
E50.6=Nimzoindiskt: 4.e3 O-O 5.Nf3 c5 6.Be2
E50.7=Nimzoindiskt: 4.e3 O-O 5.Nf3 c5 6.Bd3 Nc6
E50.8=Nimzoindiskt: 4.e3 O-O 5.Nf3 c5 6.Bd3 Nc6 7.O-O
E51.1=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5
E51.2=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.a3
E51.3=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Be2
E51.4=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Bd3
E51.5=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Bd3 Nc6
E51.6=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Bd3 Nc6 7.O-O
E51.7=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Bd3 Nc6 7.O-O a6
E51.8=Nimzoindiskt: 4.e3 O-O 5.Nf3 d5 6.Bd3 Nc6 7.O-O dxc4
E52.1=Nimzoindiskt: Huvudvarianten, 6...b6
E52.2=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O
E52.3=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7
E52.4=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.a3
E52.5=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.a3 Bd6
E52.6=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.cxd5
E52.7=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.cxd5 exd5
E52.8=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.cxd5 exd5 9.Ne5
E52.9=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.cxd5 exd5 9.a3
E52.10=Nimzoindiskt: Huvudvarianten, 6...b6 7.O-O Bb7 8.cxd5 exd5 9.a3 Bd6
E53.1=Nimzoindiskt: Huvudvarianten, 6...c5
E53.2=Nimzoindiskt: Huvudvarianten, 6...c5 7.a3
E53.3=Nimzoindiskt: Huvudvarianten, 6...c5 7.O-O
E53.4=Nimzoindiskt: Huvudvarianten, 7...Bd7
E53.5=Nimzoindiskt: Huvudvarianten, 7...Nbd7
E53.6=Nimzoindiskt: Huvudvarianten, Keresvarianten
E53.7=Nimzoindiskt: Huvudvarianten, Keres, 8.cxd5 exd5
E54.1=Nimzoindiskt: Huvudvarianten, 7...dxc4
E54.2=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4
E54.3=Nimzoindiskt: Huvudvarianten, Smyslovvarianten
E54.4=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4 Nc6
E54.5=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4 cxd4
E54.6=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4 cxd4 9.exd4
E54.7=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4 cxd4 9.exd4 a6
E54.8=Nimzoindiskt: Huvudvarianten, 7...dxc4 8.Bxc4 cxd4 9.exd4 a6 10.Bg5
E54.9=Nimzoindiskt: Huvudvarianten, Karpovvarianten
E54.10=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5
E54.11=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5 Bb7
E54.12=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5 Bb7 11.Ne5
E54.13=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5 Bb7 11.Re1
E54.14=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5 Bb7 11.Rc1
E54.15=Nimzoindiskt: Huvudvarianten, Karpov, 10.Bg5 Bb7 11.Qe2
E55.1=Nimzoindiskt: Huvudvarianten, Bronsteinvarianten
E55.2=Nimzoindiskt: Huvudvarianten, Bronstein, 9.Ne2
E55.3=Nimzoindiskt: Huvudvarianten, Bronstein, 9.a3
E55.4=Nimzoindiskt: Huvudvarianten, Bronstein, 9.a3 cd4 10.ed4
E55.5=Nimzoindiskt: Huvudvarianten, Bronstein, 9.Qe2
E55.6=Nimzoindiskt: Huvudvarianten, Bronstein, 9.Qe2 a6
E55.7=Nimzoindiskt: Huvudvarianten, Bronstein, 9.Qe2 b6
E55.8=Nimzoindiskt: Huvudvarianten, Bronstein, 9.Qe2 b6 10.Rd1
E56.1=Nimzoindiskt: Huvudvarianten, 7...Nc6
E56.2=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.cxd5
E56.3=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3
E56.4=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 Ba5
E56.5=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 Ba5 9.cxd5
E56.6=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 cxd4
E56.7=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 cxd4 9.exd4
E56.8=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 dxc4
E56.9=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 dxc4 9.Bxc4
E56.10=Nimzoindiskt: Huvudvarianten, 7...Nc6 8.a3 dxc4 9.Bxc4 Ba5
E57.1=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4
E57.2=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4
E57.3=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7
E57.4=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Be3
E57.5=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Bf4
E57.6=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Bg5
E57.7=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Qd3
E57.8=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Re1
E57.9=Nimzoindiskt: Huvudvarianten, 8...dxc4 9.Bxc4 cxd4 10.exd4 Be7 11.Re1 a6
E58.1=Nimzoindiskt: Huvudvarianten, 8...Bxc3
E58.2=Nimzoindiskt: Huvudvarianten, 8...Bxc3
E58.3=Nimzoindiskt: Huvudvarianten, 9.bxc3 b6
E58.4=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7
E58.5=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.h3
E58.6=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.Bb2
E58.7=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.Qc2
E58.8=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.cxd5
E58.9=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.cxd5 exd5 11.a4
E58.10=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.cxd5 exd5 11.a4 Re8
E58.11=Nimzoindiskt: Huvudvarianten, 9.bxc3 Qc7 10.cxd5 exd5 11.Nh4
E59.1=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4
E59.2=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4
E59.3=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7
E59.4=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.a4
E59.5=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Qe2
E59.6=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Qc2
E59.7=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bb2
E59.8=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Be2
E59.9=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bb5
E59.10=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Ba2
E59.11=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Ba2 e5
E59.12=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bd3
E59.13=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bd3 e5 12.Qc2
E59.14=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bd3 e5 12.Qc2 Re8
E59.15=Nimzoindiskt: Huvudvarianten, 9.bxc3 dxc4 10.Bxc4 Qc7 11.Bd3 e5 12.Qc2 Re8 13.de5
E60.1=King's Indian
E60.2=Kungsindiskt: Mengarinis attack
E60.3=Kungsindiskt: 3.Bg5
E60.4=Kungsindiskt: 3.d5
E60.5=Kungsindiskt: 3.d5, Danube/Adorjans gambit
E60.6=Kungsindiskt: 3.f3
E60.7=Kungsindiskt: 3.g3
E60.8=Kungsindiskt: 3.g3
E60.9=Kungsindiskt: 3.g3
E60.10=Kungsindiskt: 3.g3
E60.11=Kungsindiskt: 3.Nf3
E60.12=Kungsindiskt: 3.Nf3 d6
E60.13=Kungsindiskt: 3.Nf3 Bg7
E60.14=Kungsindiskt: b3 system
E60.15=Kungsindiskt: b3 system
E60.16=Kungsindiskt: b3 system
E60.17=Kungsindiskt: b3 system
E60.18=Kungsindiskt: b3 system
E60.19=Kungsindiskt: b3+g3 system
E60.20=Kungsindiskt: b3+g3 system
E60.21=Kungsindiskt: Fianchetto
E60.22=Kungsindiskt: Fianchetto
E60.23=Kungsindiskt: Fianchetto utan Nc3
E60.24=Kungsindiskt: Fianchetto utan Nc3
E60.25=Kungsindiskt: Fianchetto utan Nc3
E60.26=Kungsindiskt: Fianchetto, Jugoslaviskt utan Nc3
E60.27=Kungsindiskt: Fianchetto, Jugoslaviskt utan Nc3, 7.dxc5
E60.28=Kungsindiskt: Fianchetto utan Nc3, 6...c6
E60.29=Kungsindiskt: Fianchetto utan Nc3, 6...Nc6
E60.30=Kungsindiskt: Fianchetto utan Nc3, 6...Nbd7
E60.31=Kungsindiskt: Fianchetto utan Nc3, 6...Nbd7 7.Qc2
E60.32=Kungsindiskt: Fianchetto utan Nc3, 6...Nbd7 7.Qc2 e5
E60.33=Kungsindiskt: Fianchetto utan Nc3, 6...Nbd7 7.Qc2 e5 8.Rd1 Re8
E61.1=Kungsindiskt: 3.Nc3
E61.2=Kungsindiskt: 3.Nc3 c5
E61.3=Kungsindiskt: 3.Nc3 c6
E61.4=Kungsindiskt: 3.Nc3 d6
E61.5=Kungsindiskt: 3.Nc3 Bg7
E61.6=Kungsindiskt: 4.Bf4
E61.7=Kungsindiskt: 4.Bg5
E61.8=Kungsindiskt: 4.Bg5 O-O
E61.9=Kungsindiskt: 4.Bg5 O-O 5.e3 d6
E61.10=Kungsindiskt: 4.g3
E61.11=Kungsindiskt: 4.g3 d6
E61.12=Kungsindiskt: 4.g3 d6 5.Bg2
E61.13=Kungsindiskt: 4.g3 O-O
E61.14=Kungsindiskt: 4.g3 O-O 5.Bg2
E61.15=Kungsindiskt: 4.g3 O-O 5.Bg2 d6
E61.16=Kungsindiskt: Fianchetto, Flohrvarianten
E61.17=Kungsindiskt: 4.Nf3
E61.18=Kungsindiskt: 4.Nf3 d6
E61.19=Kungsindiskt: 4.Nf3 d6 5.e3
E61.20=Kungsindiskt: Smyslovs system
E61.21=Kungsindiskt: Smyslovs system
E61.22=Kungsindiskt: 4.Nf3 O-O
E61.23=Kungsindiskt: 4.Nf3 O-O 5.g3
E61.24=Kungsindiskt: 4.Nf3 O-O 5.e3
E61.25=Kungsindiskt: 4.Nf3 O-O 5.e3 d6
E61.26=Kungsindiskt: 4.Nf3 O-O 5.e3 d6 6.Be2
E61.27=Kungsindiskt: 4.Nf3 O-O 5.e3 d6 6.Be2 c5
E61.28=Kungsindiskt: 4.Nf3 O-O 5.e3 d6 6.Be2 c5
E61.29=Kungsindiskt: 4.Nf3 O-O 5.Bf4
E61.30=Kungsindiskt: 4.Nf3 O-O 5.Bf4 d6
E61.31=Kungsindiskt: 4.Nf3 d6 5.Bf4 d6 6.h3
E61.32=Kungsindiskt: 4.Nf3 d6 5.Bf4 d6 6.e3
E61.33=Kungsindiskt: Smyslovs system
E61.34=Kungsindiskt: Smyslovs system, 5...c5
E61.35=Kungsindiskt: Smyslovs system, 5...c5 6.e3
E61.36=Kungsindiskt: Smyslovs system, 5...d6
E61.37=Kungsindiskt: Smyslovs system, 6.e3
E61.38=Kungsindiskt: Smyslovs system, 6.e3 c6
E61.39=Kungsindiskt: Smyslovs system, 6.e3 c6
E61.40=Kungsindiskt: Smyslovs system, 5...O-O 6.e3 Nbd7
E61.41=Kungsindiskt: Smyslovs system, 5...O-O 6.e3 Nbd7 7.Be2
E61.42=Kungsindiskt: Smyslovs system, 5...O-O 6.e3 Nbd7 7.Be2 c6
E61.43=Kungsindiskt: Smyslovs system, 5...O-O 6.e3 Nbd7 7.Be2 c6 8.O-O
E62.1=Kungsindiskt: Fianchettovarianten
E62.2=Kungsindiskt: Fianchettovarianten
E62.3=Kungsindiskt: Fianchettovarianten
E62.4=Kungsindiskt: Fianchetto, 6...c6
E62.5=Kungsindiskt: Fianchetto, 6...c6 7.O-O
E62.6=Kungsindiskt: Fianchetto, Larsens system
E62.7=Kungsindiskt: Fianchetto, Larsens system, 8.b3
E62.8=Kungsindiskt: Fianchetto, Kavalek/Bronsteinvarianten
E62.9=Kungsindiskt: Fianchetto, Kavalek/Bronstein, 8.h3
E62.10=Kungsindiskt: Fianchetto, Kavalek/Bronstein, 8.e4
E62.11=Kungsindiskt: Fianchetto, Kavalek/Bronstein, 8.e4 Bg4
E62.12=Kungsindiskt: Fianchetto, 6...Nc6
E62.13=Kungsindiskt: Fianchetto, 6...Nc6 7.d5
E62.14=Kungsindiskt: Fianchetto, 6...Nc6 7.O-O
E62.15=Kungsindiskt: Fianchetto, 6...Nc6 7.O-O Rb8
E62.16=Kungsindiskt: Fianchetto, Spasskyvarianten
E62.17=Kungsindiskt: Fianchetto, Spassky, 8.d5
E62.18=Kungsindiskt: Fianchetto, Simaginvarianten
E62.19=Kungsindiskt: Fianchetto, Simagin, 8.d5
E62.20=Kungsindiskt: Fianchetto, Uhlmann/Szabovarianten
E62.21=Kungsindiskt: Fianchetto, Uhlmann/Szabovarianten
E62.22=Kungsindiskt: Fianchetto, Uhlmann/Szabo, 9.e4
E63.1=Kungsindiskt: Fianchetto, Pannovarianten
E63.2=Kungsindiskt: Fianchetto, Panno, 8.Re1
E63.3=Kungsindiskt: Fianchetto, Panno, 8.e4
E63.4=Kungsindiskt: Fianchetto, Panno, 8.b3
E63.5=Kungsindiskt: Fianchetto, Panno, 8.b3 Rb8
E63.6=Kungsindiskt: Fianchetto, Panno, 8.b3 Rb8 9.Bb2
E63.7=Kungsindiskt: Fianchetto, Panno, 8.b3 Rb8 9.Nd5
E63.8=Kungsindiskt: Fianchetto, Panno, 8.h3
E63.9=Kungsindiskt: Fianchetto, Panno, 8.h3 Rb8
E63.10=Kungsindiskt: Fianchetto, Panno, 8.h3 Rb8 9.Be3
E63.11=Kungsindiskt: Fianchetto, Panno, 8.h3 Rb8 9.e4
E63.12=Kungsindiskt: Fianchetto, Panno, 8.d5
E63.13=Kungsindiskt: Fianchetto, Panno, 8.d5 Na5
E64.1=Kungsindiskt: Fianchetto, Jugoslaviskt System
E64.2=Kungsindiskt: Fianchetto, Jugoslavisk, Tidigt avbyte
E64.3=Kungsindiskt: Fianchetto, Jugoslavisk, 7.d5
E64.5=Kungsindiskt: Fianchetto, Jugoslavisk, 7.d5 e6
E64.4=Kungsindiskt: Fianchetto, Jugoslavisk, 7.d5 Na6
E65.1=Kungsindiskt: Fianchetto, Jugoslavisk, 7.O-O
E65.2=Kungsindiskt: Fianchetto, Jugoslavisk, 7.O-O cxd4
E65.3=Kungsindiskt: Fianchetto, Jugoslavisk, 7.O-O Nbd7
E65.4=Kungsindiskt: Fianchetto, Jugoslavisk, 7.O-O Nc6
E65.5=Kungsindiskt: Fianchetto, Jugoslavisk, 7.O-O Nc6 8.h3
E65.6=Kungsindiskt: Fianchetto, Jugoslavisk, Avbyte
E65.7=Kungsindiskt: Fianchetto, Jugoslavisk, Avbyte, 9.Be3
E65.8=Kungsindiskt: Fianchetto, Jugoslavisk, Avbyte, 9.Bf4
E66.1=Kungsindiskt: Fianchetto, Jugoslavisk Panno
E66.2=Kungsindiskt: Fianchetto, Jugoslavisk Panno
E66.3=Kungsindiskt: Fianchetto, Jugoslavisk Panno
E66.4=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...e5
E66.5=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6
E66.6=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6 10.Rb1
E66.7=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6 10.Rb1 Rb8
E66.8=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6 10.Qc2
E66.9=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6 10.Qc2 Rb8
E66.10=Kungsindiskt: Fianchetto, Jugoslavisk Panno, 9...a6 10.Qc2 Rb8 11.b3
E66.11=Kungsindiskt: Fianchetto, Jugoslavisk Panno, Huvudvarianten
E66.12=Kungsindiskt: Fianchetto, Jugoslavisk Panno, Huvudvarianten, 12.Bb2
E66.13=Kungsindiskt: Fianchetto, Jugoslavisk Panno, Huvudvarianten, 12.Bb2 e5
E66.14=Kungsindiskt: Fianchetto, Jugoslavisk Panno, Huvudvarianten, 12.Bb2 bxc4
E67.1=Kungsindiskt: Fianchetto med 6...Nd7
E67.2=Kungsindiskt: Fianchetto med 6...Nd7 7.O-O
E67.3=Kungsindiskt: Fianchetto med 6...Nd7 7.O-O c6
E67.4=Kungsindiskt: Fianchetto, Klassiska varianten
E67.5=Kungsindiskt: Fianchetto, Klassisk, 8.d5
E67.6=Kungsindiskt: Fianchetto, Klassisk, 8.dxe5
E67.7=Kungsindiskt: Fianchetto, Klassisk, 8.b3
E67.8=Kungsindiskt: Fianchetto, Klassisk, 8.Qc2
E67.9=Kungsindiskt: Fianchetto, Klassisk, 8.Qc2 c6
E67.10=Kungsindiskt: Fianchetto, Klassisk, 8.h3
E67.11=Kungsindiskt: Fianchetto, Klassisk, 8.h3 Re8
E67.12=Kungsindiskt: Fianchetto, Klassisk, 8.h3 c6
E68.1=Kungsindiskt: Fianchetto, Klassisk, 8.e4
E68.2=Kungsindiskt: Fianchetto, Klassisk, 8.e4 Re8
E68.3=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4
E68.4=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4 9.Nxd4 Nc5
E68.5=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4 9.Nxd4 Re8
E68.6=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4 9.Nxd4 Re8 10.h3
E68.7=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4 9.Nxd4 Re8 10.h3 Nc5
E68.8=Kungsindiskt: Fianchetto, Klassisk, 8.e4 exd4 9.Nxd4 Re8 10.h3 Nc5 11.Re1 a5
E68.9=Kungsindiskt: Fianchetto, Klassisk, 8.e4 a6
E68.10=Kungsindiskt: Fianchetto, Klassisk, 8.e4 c6
E68.11=Kungsindiskt: Fianchetto, Klassisk, 8.e4 c6 9.b3
E69.1=Kungsindiskt: Fianchetto, Klassisk, 9.h3
E69.2=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qe7
E69.3=Kungsindiskt: Fianchetto, Klassisk, 9.h3 a6
E69.4=Kungsindiskt: Fianchetto, Klassisk, 9.h3 a5
E69.5=Kungsindiskt: Fianchetto, Klassisk, 9.h3 exd4
E69.6=Kungsindiskt: Fianchetto, Klassisk, 9.h3 exd4 10.Nxd4 Re8
E69.7=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qa5
E69.8=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qa5 10.Re1
E69.9=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qa5 10.Re1 exd4
E69.10=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qa5 10.Re1 exd4
E69.11=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6
E69.12=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.d5
E69.13=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.c5
E69.14=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.Re1
E69.15=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.Re1 Re8
E69.16=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.Re1 exd4
E69.17=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.Re1 exd4
E69.18=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Qb6 10.Re1 exd4 11.Nxd4 Re8
E69.19=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8
E69.20=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.b3
E69.21=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Be3
E69.22=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Be3 exd4
E69.23=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Be3 exd4 11.Nxd4
E69.24=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1
E69.25=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 Qc7
E69.26=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 a5
E69.27=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 a5 11.Be3
E69.28=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4
E69.29=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4
E69.30=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4, 11...a5
E69.31=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4, 11...Nc5
E69.32=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4, 11...Nc5 12.Rb1
E69.33=Kungsindiskt: Fianchetto, Klassisk, 9.h3 Re8 10.Re1 exd4, 11...Nc5 12.b3
E70.1=Kungsindiskt: 4.e4
E70.2=Kungsindiskt: 4.e4 O-O
E70.3=Kungsindiskt: 4.e4 O-O 5.e5
E70.4=Kungsindiskt: 4.e4 O-O 5.Nf3
E70.5=Kungsindiskt: 4.e4 d6
E70.6=Kungsindiskt: Kramer
E70.7=Kungsindiskt: Kramer, 5...O-O
E70.8=Kungsindiskt: Kramer, 5...O-O 6.Ng3
E70.9=Kungsindiskt: Kramer, 5...O-O 6.Ng3 e5
E70.10=Kungsindiskt: Kramer, 5...O-O 6.Ng3 e5 7.d5
E70.11=Kungsindiskt: 4.e4 d6 5.Bd3
E70.12=Kungsindiskt: 4.e4 d6 5.Bd3 e5
E70.13=Kungsindiskt: 4.e4 d6 5.Bd3 O-O
E70.14=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2
E70.15=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 Nc6
E70.16=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 Nc6 7.O-O
E70.17=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 Nc6 7.O-O e5
E70.18=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 c5
E70.19=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 c5 7.d5
E70.20=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 c5 7.d5 e6
E70.21=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 c5 7.d5 e6 8.O-O
E70.22=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 e5
E70.23=Kungsindiskt: 4.e4 d6 5.Bd3 O-O 6.Nge2 e5 7.d5
E70.24=Kungsindiskt: Accelererat Averbakh-system
E70.25=Kungsindiskt: Accelererat Averbakh, 5...h6
E70.26=Kungsindiskt: Accelererat Averbakh, 5...O-O
E70.27=Kungsindiskt: Accelererat Averbakh, 5...O-O 6.Qd2
E71.1=Kungsindiskt: Makagonovs system
E71.2=Kungsindiskt: Makagonov, 5...c5
E71.3=Kungsindiskt: Makagonov, 5...Nbd7
E71.4=Kungsindiskt: Makagonov, 5...O-O
E71.5=Kungsindiskt: Makagonov, 5...O-O 6.Be3
E71.6=Kungsindiskt: Makagonov, 5...O-O 6.Be3 e5
E71.7=Kungsindiskt: Makagonov, 5...O-O 6.Bg5
E71.8=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 c6
E71.9=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 h6
E71.10=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 Nbd7
E71.11=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 Na6
E71.12=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 Na6 7.Bd3
E71.13=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 Na6 7.Bd3 e5
E71.14=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 c5
E71.15=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 c5 7.d5
E71.16=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 c5 7.d5 b5
E71.17=Kungsindiskt: Makagonov, 5...O-O 6.Bg5 c5 7.d5 e6
E72.1=Kungsindiskt: 4.e4 d6 5.g3
E72.2=Kungsindiskt: 4.e4 d6 5.g3 O-O
E72.3=Kungsindiskt: 4.e4 d6 5.g3 O-O 6.Bg2
E72.4=Kungsindiskt: 4.e4 d6 5.g3 O-O 6.Bg2 Nbd7
E72.5=Kungsindiskt: 4.e4 d6 5.g3 O-O 6.Bg2 Nc6
E72.6=Kungsindiskt: 4.e4 d6 5.g3 O-O 6.Bg2 c5
E72.7=Kungsindiskt: 4.e4 d6 5.g3 O-O 6.Bg2 e5
E72.8=Kungsindiskt: Pomarsystemet
E72.9=Kungsindiskt: Pomarsystemet
E73.1=Kungsindiskt: 5.Be2
E73.2=Kungsindiskt: 5.Be2 c5
E73.3=Kungsindiskt: 5.Be2 e5
E73.4=Kungsindiskt: 5.Be2 e5 6.d5
E73.5=Kungsindiskt: 5.Be2 Nbd7
E73.6=Kungsindiskt: 5.Be2 O-O
E73.7=Kungsindiskt: 5.Be2 O-O 6.g4
E73.8=Kungsindiskt: Semi-Averbakhsystemet
E73.9=Kungsindiskt: Averbakh
E73.10=Kungsindiskt: Averbakh, 6...c6
E73.11=Kungsindiskt: Averbakh, 6...c6 7.Qd2
E73.12=Kungsindiskt: Averbakh, 6...c6 7.Qd2 Nbd7
E73.13=Kungsindiskt: Averbakh, 6...Nbd7
E73.14=Kungsindiskt: Averbakh, 6...Nbd7 7.Qd2
E73.15=Kungsindiskt: Averbakh, 6...Nbd7 7.Qd2 e5
E73.16=Kungsindiskt: Averbakh, 6...Nbd7 7.Qd2 e5 8.d5
E73.17=Kungsindiskt: Averbakh, 6...Nbd7 7.Qd2 e5 8.d5 Nc5
E73.18=Kungsindiskt: Averbakh, 6...Na6
E73.19=Kungsindiskt: Averbakh, 6...Na6 7.h4
E73.20=Kungsindiskt: Averbakh, 6...Na6 7.Qd2
E73.21=Kungsindiskt: Averbakh, 6...Na6 7.Qd2 e5
E73.22=Kungsindiskt: Averbakh, 6...Na6 7.Qd2 e5 8.d5
E73.23=Kungsindiskt: Averbakh, 6...Na6 7.Qd2 e5 8.d5 c6
E73.24=Kungsindiskt: Averbakh, 6...Na6 7.Qd2 e5 8.d5 Qe8
E73.25=Kungsindiskt: Averbakh, 6...h6
E73.26=Kungsindiskt: Averbakh, 6...h6 7.Be3
E73.27=Kungsindiskt: Averbakh, 6...h6 7.Be3 c5
E73.28=Kungsindiskt: Averbakh, 6...h6 7.Be3 e5
E73.29=Kungsindiskt: Averbakh, 6...h6 7.Be3 e5 8.d5
E73.30=Kungsindiskt: Averbakh, 6...h6 7.Be3 e5 8.d5 c6
E73.31=Kungsindiskt: Averbakh, 6...h6 7.Be3 e5 8.d5 Nbd7
E74.1=Kungsindiskt: Averbakh, 6...c5
E74.2=Kungsindiskt: Averbakh, 6...c5 7.dxc5
E74.3=Kungsindiskt: Averbakh, 6...c5 7.dxc5 Qa5
E74.4=Kungsindiskt: Averbakh, 6...c5 7.dxc5 Qa5 8.Bd2 Qxc5 9.Nf3 Bg4
E74.5=Kungsindiskt: Averbakh, 6...c5 7.d5
E74.6=Kungsindiskt: Averbakh, 6...c5 7.d5 Qa5
E74.7=Kungsindiskt: Averbakh, 6...c5 7.d5 b5
E74.8=Kungsindiskt: Averbakh, 6...c5 7.d5 b5 8.cxb5 a6 9.a4
E74.9=Kungsindiskt: Averbakh, 6...c5 7.d5 a6
E74.10=Kungsindiskt: Averbakh, 6...c5 7.d5 a6 8.a4
E74.11=Kungsindiskt: Averbakh, 6...c5 7.d5 a6 8.a4 Qa5
E74.12=Kungsindiskt: Averbakh, 6...c5 7.d5 h6
E74.13=Kungsindiskt: Averbakh, 6...c5 7.d5 h6 8.Bh4
E74.14=Kungsindiskt: Averbakh, 6...c5 7.d5 h6 8.Be3
E74.15=Kungsindiskt: Averbakh, 6...c5 7.d5 h6 8.Be3 e6
E74.16=Kungsindiskt: Averbakh, 6...c5 7.d5 h6 8.Bf4
E74.17=Kungsindiskt: Averbakh, 6...c5 7.d5 h6 8.Bf4 e6
E75.1=Kungsindiskt: Averbakh, 7.d5 e6
E75.2=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3
E75.3=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 exd5
E75.4=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 exd5 9.exd5
E75.5=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 h6
E75.6=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 h6 9.Bd2
E75.7=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 h6 9.Be3
E75.8=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 h6 9.Bf4
E75.9=Kungsindiskt: Averbakh, 7.d5 e6 8.Nf3 h6 9.Bh4
E75.10=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2
E75.11=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5
E75.12=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5 9.exd5
E75.13=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5 9.exd5 a6
E75.14=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5 9.exd5 Re8
E75.15=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5 9.exd5 Re8 10.Nf3
E75.16=Kungsindiskt: Averbakh, 7.d5 e6 8.Qd2 exd5 9.exd5 Re8 10.Nf3 Bg4
E76.1=Kungsindiskt: Fyrbondeattack
E76.2=Kungsindiskt: Fyrbondeattack, 5...c5
E76.3=Kungsindiskt: Fyrbondeattack, Avbyte
E76.4=Kungsindiskt: Fyrbondeattack, 5...c5 6.d5
E76.5=Kungsindiskt: Fyrbondeattack, 5...O-O
E76.6=Kungsindiskt: Fyrbondeattack, 5...O-O 6.Nf3
E76.7=Kungsindiskt: Fyrbondeattack, 6.Nf3 Bg4
E76.8=Kungsindiskt: Fyrbondeattack, 6.Nf3 Na6
E76.9=Kungsindiskt: Fyrbondeattack, 6.Nf3 Na6 7.e5
E76.10=Kungsindiskt: Fyrbondeattack, 6.Nf3 Na6 7.Be2
E76.11=Kungsindiskt: Fyrbondeattack, 6.Nf3 Na6 7.Bd3
E76.12=Kungsindiskt: Fyrbondeattack, 6.Nf3 Na6 7.Bd3 e5
E76.13=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5
E76.14=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.dxc5
E76.15=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.dxc5 Qa5 8.Bd3 Qxc5 9.Qe2 Nc6
E76.16=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5
E76.17=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5 a6
E76.18=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5 b5
E76.19=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5 b5 8.cxb5 a6 9.a4
E76.20=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5 e6
E76.21=Kungsindiskt: Fyrbondeattack, 6.Nf3 c5 7.d5 e6 8.dxe6
E77.1=Kungsindiskt: Fyrbondeattack, 6.Be2
E77.2=Kungsindiskt: Fyrbondeattack, 6.Be2 c5
E77.3=Kungsindiskt: Fyrbondeattack, 6.Be2 c5 7.d5
E77.4=Kungsindiskt: Fyrbondeattack, Sexbonde-varianten
E77.5=Kungsindiskt: Fyrbondeattack, 6.Be2 c5 7.d5 e6 8.Nf3
E77.6=Kungsindiskt: Fyrbondeattack, 6.Be2 c5 7.d5 e6 8.Nf3 exd5 9.exd5
E77.7=Kungsindiskt: Fyrbondeattack, Florentines gambit
E78.1=Kungsindiskt: Fyrbondeattack, 7.Nf3
E78.2=Kungsindiskt: Fyrbondeattack, 7.Nf3 Bg4
E78.3=Kungsindiskt: Fyrbondeattack, 7.Nf3 cxd4
E78.4=Kungsindiskt: Fyrbondeattack, 7.Nf3 cxd4
E79.1=Kungsindiskt: Fyrbondeattack, Huvudvarianten
E79.2=Kungsindiskt: Fyrbondeattack, Huvudvarianten, 9...Nxd4
E79.3=Kungsindiskt: Fyrbondeattack, Huvudvarianten, 9...Bd7
E79.4=Kungsindiskt: Fyrbondeattack, Huvudvarianten, 9...Bd7 10.Qd2
E80.1=Kungsindiskt: S�mischvarianten
E80.2=Kungsindiskt: S�misch, 5...Na6
E80.3=Kungsindiskt: S�misch, 5...Nc6
E80.4=Kungsindiskt: S�misch, 5...Nbd7
E80.5=Kungsindiskt: S�misch, 5...e5
E80.6=Kungsindiskt: S�misch, 5...e5 6.Nge2
E80.7=Kungsindiskt: S�misch, 5...e5 6.d5
E80.8=Kungsindiskt: S�misch, 5...c5
E80.9=Kungsindiskt: S�misch, 5...c5 Dambyte
E80.10=Kungsindiskt: S�misch, 5...a6
E80.11=Kungsindiskt: S�misch, 5...a6 6.Be3
E80.12=Kungsindiskt: S�misch, 5...c6
E80.13=Kungsindiskt: S�misch, 5...c6 6.Be3
E80.14=Kungsindiskt: S�misch, 5...c6 6.Be3 a6
E80.15=Kungsindiskt: S�misch, 5...c6 6.Be3 a6 7.a4
E80.16=Kungsindiskt: S�misch, 5...c6 6.Be3 a6 7.Bd3
E81.1=Kungsindiskt: S�misch, 5...O-O
E81.2=Kungsindiskt: S�misch, 5...O-O 6.Nge2
E81.3=Kungsindiskt: S�misch, 5...O-O 6.Nge2 e5
E81.4=Kungsindiskt: S�misch, 5...O-O 6.Nge2 c5
E81.5=Kungsindiskt: S�misch, 5...O-O 6.Nge2 c5 7.d5
E81.6=Kungsindiskt: S�misch, 5...O-O 6.Bg5
E81.7=Kungsindiskt: S�misch, 5...O-O 6.Bg5 Nc6
E81.8=Kungsindiskt: S�misch, 5...O-O 6.Bg5 a6
E81.9=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5
E81.10=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5 7.d5
E81.11=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5 7.d5 a6
E81.12=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5 7.d5 h6
E81.13=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5 7.d5 e6
E81.14=Kungsindiskt: S�misch, 5...O-O 6.Bg5 c5 7.d5 e6 8.Qd2
E81.15=Kungsindiskt: S�misch, 5...O-O 6.Be3
E81.16=Kungsindiskt: S�misch, 5...O-O 6.Be3 a6
E81.17=Kungsindiskt: S�misch, 5...O-O 6.Be3 a6 7.Qd2
E81.18=Kungsindiskt: S�misch, 5...O-O 6.Be3 c6
E81.19=Kungsindiskt: S�misch, Byrnevarianten
E81.20=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5
E81.21=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 7.d5
E81.22=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 7.dxc5
E81.23=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 Dambyte
E81.24=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 7.Nge2
E81.25=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 7.Nge2 Nc6
E81.26=Kungsindiskt: S�misch, 5...O-O 6.Be3 c5 7.Nge2 Nc6 8.d5
E81.27=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7
E81.28=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7 7.Qd2
E81.29=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7 7.Qd2 c5
E81.30=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7 7.Qd2 c5 8.d5
E81.31=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7 7.Qd2 c5 8.Nge2
E81.32=Kungsindiskt: S�misch, 5...O-O 6.Be3 Nbd7 7.Qd2 c5 8.Nge2 a6
E82.1=Kungsindiskt: S�misch, Fianchetto
E82.2=Kungsindiskt: S�misch, Fianchetto, 7.Qd2
E82.3=Kungsindiskt: S�misch, Fianchetto, Bronsteinvarianten
E82.4=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 Bb7
E82.5=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 Bb7 8.Nge2 c5
E82.6=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 Bb7 8.Nge2 c5 9.d5 e6
E82.8=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 a6
E82.9=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 a6 8.Nge2 c5
E82.11=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 a6 8.Nge2 c5 9.d5
E82.10=Kungsindiskt: S�misch, Fianchetto, 7.Bd3 a6 8.Nge2 c5 9.e5
E83.1=Kungsindiskt: S�misch, 6...Nc6
E83.2=Kungsindiskt: S�misch, 6...Nc6 7.Qd2
E83.3=Kungsindiskt: S�misch, 6...Nc6 7.Qd2 a6 8.O-O-O
E83.4=Kungsindiskt: S�misch, 6...Nc6 7.Nge2
E83.5=Kungsindiskt: S�misch, Rubanvarianten
E83.6=Kungsindiskt: S�misch, Ruban, 8.Qd2 Re8
E83.7=Kungsindiskt: S�misch, Panno
E83.8=Kungsindiskt: S�misch, Panno, 8.a3
E83.9=Kungsindiskt: S�misch, Panno, 8.Nc1
E83.10=Kungsindiskt: S�misch, Panno, 8.Qd2
E84.1=Kungsindiskt: S�misch, Panno Huvudvarianten
E84.2=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.O-O-O
E84.3=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Rb1
E84.4=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Bh6
E84.5=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Nc1
E84.6=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Nc1 e5
E84.7=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Nc1 e5 10.Nb3
E84.8=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.Nc1 e5 10.d5
E84.9=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.h4
E84.10=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.h4 b5
E84.11=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.h4 h5
E84.12=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.h4 h5 10.O-O-O
E84.13=Kungsindiskt: S�misch, Panno Huvudvarianten, 9.h4 h5 10.O-O-O b5 11.Bh6
E85.1=Kungsindiskt: S�misch, Orthodoxvarianten
E85.2=Kungsindiskt: S�misch, Orthodox, 7.dxe5
E85.3=Kungsindiskt: S�misch, Orthodox, Dambyte
E85.4=Kungsindiskt: S�misch, Orthodox, 7.Nge2
E85.5=Kungsindiskt: S�misch, Orthodox, 7.Nge2 exd4
E85.6=Kungsindiskt: S�misch, Orthodox, 7.Nge2 Nbd7
E85.7=Kungsindiskt: S�misch, Orthodox, 7.Nge2 Nc6
E85.8=Kungsindiskt: S�misch, Orthodox, 7.Nge2 Nc6 8.d5
E86.1=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6
E86.2=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.d5
E86.3=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qb3
E86.4=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2
E86.5=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2 Nbd7
E86.6=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2 Nbd7 9.d5
E86.7=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2 Nbd7 9.O-O-O
E86.8=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2 Nbd7 9.O-O-O a6
E86.9=Kungsindiskt: S�misch, Orthodox, 7.Nge2 c6 8.Qd2 Nbd7 9.O-O-O a6 10.Kb1
E87.1=Kungsindiskt: S�misch, Orthodox, 7.d5
E87.2=Kungsindiskt: S�misch, Orthodox, 7.d5 a5
E87.3=Kungsindiskt: S�misch, Orthodox, 7.d5 Nbd7
E87.4=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5
E87.5=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5 8.Qd2
E87.6=Kungsindiskt: S�misch, Orthodox, Bronsteinvarianten
E87.7=Kungsindiskt: S�misch, Orthodox, Bronstein, 9.g3
E87.8=Kungsindiskt: S�misch, Orthodox, Bronstein, 9.Bf2
E87.9=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5 8.Qd2 f5
E87.10=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5 8.Qd2 f5 9.O-O-O
E87.11=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5 8.Qd2 f5 9.O-O-O f4
E87.12=Kungsindiskt: S�misch, Orthodox, 7.d5 Nh5 8.Qd2 f5 9.O-O-O Nd7
E88.1=Kungsindiskt: S�misch, Orthodox, 7.d5 c6
E88.6=Kungsindiskt: S�misch, Orthodox, 7.d5 c6 8.Qd2
E88.7=Kungsindiskt: S�misch, Orthodox, 7.d5 c6 8.Qd2 cxd5
E88.8=Kungsindiskt: S�misch, Orthodox, 7.d5 c6 8.Qd2 cxd5 9.cxd5 a6
E88.9=Kungsindiskt: S�misch, Orthodox, 7.d5 c6 8.Qd2 cxd5 9.cxd5 a6 10.Bd3
E88.2=Kungsindiskt: S�misch, Orthodox, Polugayevsky
E88.3=Kungsindiskt: S�misch, Orthodox, Polugayevsky, 8...b5
E88.4=Kungsindiskt: S�misch, Orthodox, Polugayevsky, 8...cxd5
E88.5=Kungsindiskt: S�misch, Orthodox, Polugayevsky, 8...cxd5 9.cxd5 Nh5
E89.1=Kungsindiskt: S�misch, Orthodox Huvudvarianten
E89.2=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 9...a6
E89.3=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 9...Bd7
E89.4=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 9...Nbd7
E89.5=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 10.Qd2
E89.6=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 10.Qd2 a6
E89.7=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 10.Qd2 a6 11.g4
E89.8=Kungsindiskt: S�misch, Orthodox Huvudvarianten, 10.Qd2 a6 11.g4 h5
E90.1=Kungsindiskt: 5.Nf3
E90.2=Kungsindiskt: 5.Nf3 Nbd7
E90.3=Kungsindiskt: 5.Nf3 Nbd7 6.Be2
E90.4=Kungsindiskt: 5.Nf3 Nbd7 6.Be2 e5
E90.5=Kungsindiskt: 5.Nf3 Bg4
E90.6=Kungsindiskt: 5.Nf3 c5
E90.7=Kungsindiskt: 5.Nf3 c5 6.d5 O-O
E90.8=Kungsindiskt: 5.Nf3 O-O
E90.9=Kungsindiskt: 5.Nf3 O-O 6.Bd3
E90.10=Kungsindiskt: Zinnowitzvarianten
E90.11=Kungsindiskt: Zinnowitz, 6...h6
E90.12=Kungsindiskt: Larsenvarianten
E90.13=Kungsindiskt: Larsen, 6...c5
E90.14=Kungsindiskt: Larsen, 6...e5
E90.15=Kungsindiskt: Larsen, 6...e5, Dambyte
E90.16=Kungsindiskt: 5.Nf3 O-O 6.h3
E90.17=Kungsindiskt: 5.Nf3 O-O 6.h3 Nbd7
E90.18=Kungsindiskt: 5.Nf3 O-O 6.h3 Nbd7 7.Bg5
E90.19=Kungsindiskt: 5.Nf3 O-O 6.h3 Na6
E90.20=Kungsindiskt: 5.Nf3 O-O 6.h3 Na6 7.Bg5
E90.21=Kungsindiskt: 5.Nf3 O-O 6.h3 e5
E90.22=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.Be3
E90.23=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 Dambyte
E90.24=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5
E90.25=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 a5
E90.26=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Nbd7
E90.27=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Nbd7 8.Be3
E90.28=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Nbd7 8.Bg5
E90.29=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Na6
E90.30=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Na6 8.Be3
E90.31=Kungsindiskt: 5.Nf3 O-O 6.h3 e5 7.d5 Na6 8.Bg5
E90.32=Kungsindiskt: 5.Nf3 O-O 6.h3 c5
E90.33=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.Be3
E90.34=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5
E90.35=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6
E90.36=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3
E90.37=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 Na6
E90.38=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 Na6 9.O-O
E90.39=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 Na6 9.O-O Nc7
E90.40=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 exd5
E90.41=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 exd5 9.exd5
E90.42=Kungsindiskt: 5.Nf3 O-O 6.h3 c5 7.d5 e6 8.Bd3 exd5 9.exd5 Re8
E91.1=Kungsindiskt: 6.Be2
E91.2=Kungsindiskt: 6.Be2 a5
E91.3=Kungsindiskt: 6.Be2 a6
E91.4=Kungsindiskt: 6.Be2 c6
E91.5=Kungsindiskt: 6.Be2 c6 7.O-O
E91.6=Kungsindiskt: 6.Be2 c5
E91.7=Kungsindiskt: 6.Be2 c5 7.d5
E91.8=Kungsindiskt: 6.Be2 c5 7.d5 e6
E91.9=Kungsindiskt: 6.Be2 c5 7.d5 e6 8.O-O
E91.10=Kungsindiskt: 6.Be2 c5 7.d5 e6 8.O-O Re8
E91.11=Kungsindiskt: 6.Be2 c5 7.d5 e6 8.O-O Re8 9.Nd2
E91.12=Kungsindiskt: 6.Be2 c5 7.O-O
E91.13=Kungsindiskt: 6.Be2 c5 7.O-O Nc6
E91.14=Kungsindiskt: Kasackvarianten
E91.15=Kungsindiskt: Kasackvarianten, 7.Bg5
E91.16=Kungsindiskt: Kasackvarianten, 7.O-O
E91.17=Kungsindiskt: Kasackvarianten, 7.O-O c5
E91.18=Kungsindiskt: Kasackvarianten, 7.O-O c6
E91.19=Kungsindiskt: 6.Be2 Nc6
E91.20=Kungsindiskt: 6.Be2 Nc6 7.d5
E91.21=Kungsindiskt: 6.Be2 Nbd7
E91.22=Kungsindiskt: 6.Be2 Nbd7 7.Bg5
E91.23=Kungsindiskt: 6.Be2 Nbd7 7.e5
E91.24=Kungsindiskt: 6.Be2 Nbd7 7.O-O
E91.25=Kungsindiskt: 6.Be2 Nbd7 7.O-O c6
E91.26=Kungsindiskt: 6.Be2 Bg4
E91.27=Kungsindiskt: 6.Be2 Bg4 7.Be3
E91.28=Kungsindiskt: 6.Be2 Bg4 7.Be3 Nfd7
E91.29=Kungsindiskt: 6.Be2 Bg4 7.Be3 Nfd7 8.Rc1
E91.30=Kungsindiskt: 6.Be2 Bg4 7.Be3 Nfd7 8.Ng1
E92.1=Kungsindiskt: 6.Be2 e5
E92.2=Kungsindiskt: 6.Be2 e5 Dambyte
E92.3=Kungsindiskt: 6.Be2 e5 Dambyte
E92.4=Kungsindiskt: 6.Be2 e5 Dambyte, 9.Bg5
E92.5=Kungsindiskt: 6.Be2 e5 Dambyte, 9.Bg5 c6
E92.6=Kungsindiskt: 6.Be2 e5 Dambyte, 9.Bg5 Re8
E92.7=Kungsindiskt: 6.Be2 e5 Dambyte, 9.Bg5 Re8 10.Nd5
E92.8=Kungsindiskt: Gligoric-Taimanov-systemet
E92.9=Kungsindiskt: Gligoric-Taimanov, 7...c6
E92.10=Kungsindiskt: Gligoric-Taimanov, 7...exd4
E92.11=Kungsindiskt: Gligoric-Taimanov, 7...Qe7
E92.12=Kungsindiskt: Gligoric-Taimanov, 7...Ng4
E92.13=Kungsindiskt: Gligoric-Taimanov, 7...Ng4 8.Bg5 f6 9.Bc1
E92.14=Kungsindiskt: Gligoric-Taimanov, 7...Ng4 8.Bg5 f6 9.Bh4
E92.15=Kungsindiskt: Gligoric-Taimanov, Huvudvarianten
E92.16=Kungsindiskt: Petrosians system
E92.17=Kungsindiskt: Petrosian, 7...c5
E92.18=Kungsindiskt: Petrosian, 7...c5 8.Bg5
E92.19=Kungsindiskt: Petrosian, Steinvarianten
E92.20=Kungsindiskt: Petrosian, Stein, 8.h3
E92.21=Kungsindiskt: Petrosian, Stein, 8.Bg5
E92.22=Kungsindiskt: Petrosian, Stein, 8.Bg5 h6
E92.23=Kungsindiskt: Petrosian, Stein, 8.Bg5 h6 9.Bh4 Na6
E92.24=Kungsindiskt: Petrosian, Stein, Huvudvarianten
E92.25=Kungsindiskt: Petrosian, Stein, Huvudvarianten, 10...Qe8
E92.26=Kungsindiskt: Petrosian, Stein, Huvudvarianten, 10...Qe8 11.O-O
E92.27=Kungsindiskt: Petrosian, Stein, Huvudvarianten, 10...Qe8 11.O-O Bd7
E92.28=Kungsindiskt: Petrosian, Stein, Huvudvarianten, 10...Qe8 11.O-O Nh7
E93.1=Kungsindiskt: Petrosian, Huvudvarianten
E93.2=Kungsindiskt: Petrosian, Huvudvarianten, 8.Qc2
E93.3=Kungsindiskt: Petrosian, Huvudvarianten, 8.Be3
E93.4=Kungsindiskt: Petrosian, Huvudvarianten, 8.Be3 Ng4
E93.5=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5
E93.6=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5 h6
E93.7=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5 h6 9.Bh4
E93.8=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5 h6 9.Bh4 a6
E93.9=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5 h6 9.Bh4 a5
E93.10=Kungsindiskt: Petrosian, Huvudvarianten, 8.Bg5 h6 9.Bh4 g5
E93.11=Kungsindiskt: Petrosian, Keresvarianten
E94.1=Kungsindiskt: 7.O-O
E94.2=Kungsindiskt: 7.O-O exd4
E94.3=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3
E94.4=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3 c6
E94.5=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3 c6 10.Kh1
E94.6=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3 Nc6
E94.7=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3 Nc6 10.Be3
E94.8=Kungsindiskt: 7.O-O exd4 8.Nxd4 Re8 9.f3 Nc6 10.Be3 Nh5 11.Qd2
E94.9=Kungsindiskt: Donnervarianten
E94.10=Kungsindiskt: Donner, 8.d5
E94.11=Kungsindiskt: Donner, 8.Be3
E94.12=Kungsindiskt: Glekvarianten
E94.13=Kungsindiskt: Glek, 8.Re1
E94.14=Kungsindiskt: Glek, 8.Re1 c6
E94.15=Kungsindiskt: Glek, 8.Re1 c6 9.Bf1
E94.16=Kungsindiskt: Glek, 8.Be3
E94.17=Kungsindiskt: Glek, 8.Be3 Ng4
E94.18=Kungsindiskt: Glek, 8.Be3 Ng4 9.Ng5 Qe8
E94.19=Kungsindiskt: Glek, Huvudvarianten
E94.20=Kungsindiskt: Glek, Huvudvarianten, 11.h3
E94.21=Kungsindiskt: Glek, Huvudvarianten, 11.h3 h6
E94.22=Kungsindiskt: 7.O-O Nbd7
E94.23=Kungsindiskt: 7.O-O Nbd7 8.d5
E94.24=Kungsindiskt: 7.O-O Nbd7 8.d5 Nc5
E94.25=Kungsindiskt: 7.O-O Nbd7 8.d5 Nc5 9.Qc2
E94.26=Kungsindiskt: 7.O-O Nbd7 8.d5 Nc5 9.Qc2 a5
E94.27=Kungsindiskt: 7.O-O Nbd7 8.Qc2
E94.28=Kungsindiskt: 7.O-O Nbd7 8.Qc2 Re8
E94.29=Kungsindiskt: 7.O-O Nbd7 8.Qc2 c6
E94.30=Kungsindiskt: 7.O-O Nbd7 8.Be3
E94.31=Kungsindiskt: 7.O-O Nbd7 8.Be3 Ng4
E94.32=Kungsindiskt: 7.O-O Nbd7 8.Be3 Re8
E94.33=Kungsindiskt: 7.O-O Nbd7 8.Be3 c6
E94.34=Kungsindiskt: 7.O-O Nbd7 8.Be3 c6 9.d5
E94.35=Kungsindiskt: 7.O-O Nbd7 8.Be3 c6 9.d5 c5
E95.1=Kungsindiskt: 7.O-O Nbd7 8.Re1
E95.2=Kungsindiskt: 7.O-O Nbd7 8.Re1 a5
E95.3=Kungsindiskt: 7.O-O Nbd7 8.Re1 h6
E95.4=Kungsindiskt: 7.O-O Nbd7 8.Re1 Re8
E95.5=Kungsindiskt: 7.O-O Nbd7 8.Re1 Re8 9.Bf1
E95.6=Kungsindiskt: 7.O-O Nbd7 8.Re1 exd4
E95.7=Kungsindiskt: 7.O-O Nbd7 8.Re1 exd4 9.Nxd4 Nc5
E95.8=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6
E95.9=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Rb1
E95.10=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Bf1
E95.11=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Bf1 Re8
E95.12=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Bf1 exd4
E95.13=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Bf1 exd4 10.Nxd4 Ng4
E95.14=Kungsindiskt: 7.O-O Nbd7 8.Re1 c6 9.Bf1 exd4 10.Nxd4 Re8
E96.1=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten
E96.2=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.h3
E96.3=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.dxe5
E96.4=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.dxe5
E96.5=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.Rb1
E96.6=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.Rb1 Re8
E96.7=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.Rb1 Re8 11.d5
E96.8=Kungsindiskt: 7.O-O Nbd7, Gamla huvudvarianten, 10.Rb1 Re8 11.d5 Nc5 12.b3
E97.1=Kungsindiskt: Mar del Plata
E97.2=Kungsindiskt: Mar del Plata, 8.dxe5
E97.3=Kungsindiskt: Mar del Plata, 8.Be3
E97.4=Kungsindiskt: Mar del Plata, 8.Be3 Ng4
E97.5=Kungsindiskt: Mar del Plata, 8.Be3 Ng4
E97.6=Kungsindiskt: Mar del Plata, 8.d5
E97.7=Kungsindiskt: Mar del Plata, 8.d5 Ne7
E97.8=Kungsindiskt: Mar del Plata, Odessavarianten
E97.9=Kungsindiskt: Mar del Plata, 9.Bd2
E97.10=Kungsindiskt: Mar del Plata, Barjonettattack
E97.11=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Kh8
E97.12=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Ne8
E97.13=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Ne8 10.c5
E97.14=Kungsindiskt: Mar del Plata, Barjonettattack, 9...a5
E97.15=Kungsindiskt: Mar del Plata, Barjonettattack, 9...a5 10.bxa5
E97.16=Kungsindiskt: Mar del Plata, Barjonettattack, 9...a5 10.Ba3
E97.17=Kungsindiskt: Mar del Plata, Barjonettattack, 9...a5 10.Ba3 axb4
E97.18=Kungsindiskt: Mar del Plata, Barjonettattack, 9...a5 10.Ba3 axb4 11.Bxb4 Nd7
E97.19=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Nh5
E97.20=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Nh5 10.c5
E97.21=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Nh5 10.g3
E97.22=Kungsindiskt: Mar del Plata, Barjonettattack, 9...Nh5 10.Re1
E97.23=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 a5
E97.24=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 Nf4
E97.25=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 Nf4 11.Bf1 a5
E97.26=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 Nf4 11.Bf1 a5 12.bxa5
E97.27=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 f5
E97.28=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 f5 11.Ng5 Nf6
E97.29=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 f5 11.Ng5 Nf6 12.Bf3
E97.30=Kungsindiskt: Mar del Plata, Barjonett, 9...Nh5 10.Re1 f5 11.Ng5 Nf6 12.Bf3 c6
E97.31=Kungsindiskt: Mar del Plata, 9.Nd2
E97.32=Kungsindiskt: Mar del Plata, 9.Nd2 Ne8
E97.33=Kungsindiskt: Mar del Plata, 9.Nd2 Ne8 10.b4
E97.34=Kungsindiskt: Mar del Plata, 9.Nd2 Nd7
E97.35=Kungsindiskt: Mar del Plata, 9.Nd2 Nd7 10.b4
E97.36=Kungsindiskt: Mar del Plata, 9.Nd2 c5
E97.37=Kungsindiskt: Mar del Plata, 9.Nd2 a5
E97.38=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.Rb1
E97.39=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.a3
E97.40=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.a3 Bd7
E97.41=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.a3 Nd7
E97.42=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.a3 Nd7 11.Rb1
E97.43=Kungsindiskt: Mar del Plata, 9.Nd2 a5 10.a3 Nd7 11.Rb1 f5 12.b4
E98.1=Kungsindiskt: Mar del Plata, 9.Ne1
E98.2=Kungsindiskt: Mar del Plata, 9.Ne1 c5
E98.3=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8
E98.4=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8 10.Nd3
E98.5=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8 10.Nd3 f5
E98.6=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8 10.Be3
E98.7=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8 10.Be3 f5 11.f3
E98.8=Kungsindiskt: Mar del Plata, 9.Ne1 Ne8 10.Be3 f5 11.f3 f4
E98.9=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7
E98.10=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Kh1
E98.11=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Be3
E98.12=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Be3 f5
E98.13=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Nd3
E98.14=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Nd3 f5
E98.15=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Nd3 f5 11.Bd2
E98.16=Kungsindiskt: Mar del Plata, Fischervarianten
E98.17=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Nd3 f5 11.Bd2 Kh8
E98.18=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.Nd3 f5 11.Bd2 Nf6
E98.19=Kungsindiskt: Mar del Plata, 9.Ne1 Nd7 10.f3
E99.1=Kungsindiskt: Mar del Plata, 10.f3 f5
E99.2=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3
E99.3=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3 Nf6
E99.4=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3 Nf6 12.Bd2
E99.5=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3 Nf6 12.Bd2 f4
E99.6=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3 Nf6 12.Bd2 f4 13.c5
E99.7=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Nd3 f4
E99.8=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Be3
E99.9=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Be3 f4
E99.10=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Be3 f4 12.Bf2 g5
E99.11=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Be3 f4 12.Bf2 g5 13.a4
E99.12=Kungsindiskt: Mar del Plata, 10.f3 f5 11.Be3 f4 12.Bf2 g5 13.a4 Ng6
E99.13=Kungsindiskt: Mar del Plata, Benkoattack
E99.14=Kungsindiskt: Mar del Plata, Benkoattack, 11...Kh8
E99.15=Kungsindiskt: Mar del Plata, Benkoattack, 11...Nf6
E99.16=Kungsindiskt: Mar del Plata, Benkoattack, 11...Nf6 12.Nd3
